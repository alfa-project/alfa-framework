/*
 * Copyright 2025 ALFA Project. All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`timescale 1ns / 1ps

module alib_atan (
    input  signed [15:0] y,
    input  signed [15:0] x,
    output wire   [15:0] arctan_angle
);

  // Define LUT parameters
  parameter ANGLE_RANGE = 36000;  // Range of angles in tenths of degrees (-π/2 to π/2)
  parameter LUT_SIZE = 2048;  // Size of the LUT

  // Calculate y/x ratio
  wire signed [15:0] y_over_x = (x != 0) ? (y << 1) / x : (y < 0) ? -32768 : 32767;

  // Calculate index for LUT
  wire        [ 9:0] lut_index = (y_over_x < 0) ? -y_over_x : y_over_x;

  // LUT for arctangent values
  wire signed [15:0] value                                                         [LUT_SIZE - 1:0];

  // Assign output based on LUT

  assign arctan_angle = (x==0) ? (y>=0) ? 90 * (ANGLE_RANGE / 360) : 
                                         -90 * (ANGLE_RANGE / 360) :
                        (x>0) ? value[lut_index] :
                         -value[lut_index];

  initial begin

    value[0] = 15'd4500;
    value[1] = -15'd4497;
    value[2] = -15'd4494;
    value[3] = -15'd4492;
    value[4] = -15'd4489;
    value[5] = -15'd4486;
    value[6] = -15'd4483;
    value[7] = -15'd4480;
    value[8] = -15'd4478;
    value[9] = -15'd4475;
    value[10] = -15'd4472;
    value[11] = -15'd4469;
    value[12] = -15'd4466;
    value[13] = -15'd4463;
    value[14] = -15'd4461;
    value[15] = -15'd4458;
    value[16] = -15'd4455;
    value[17] = -15'd4452;
    value[18] = -15'd4449;
    value[19] = -15'd4446;
    value[20] = -15'd4443;
    value[21] = -15'd4441;
    value[22] = -15'd4438;
    value[23] = -15'd4435;
    value[24] = -15'd4432;
    value[25] = -15'd4429;
    value[26] = -15'd4426;
    value[27] = -15'd4423;
    value[28] = -15'd4421;
    value[29] = -15'd4418;
    value[30] = -15'd4415;
    value[31] = -15'd4412;
    value[32] = -15'd4409;
    value[33] = -15'd4406;
    value[34] = -15'd4403;
    value[35] = -15'd4400;
    value[36] = -15'd4397;
    value[37] = -15'd4395;
    value[38] = -15'd4392;
    value[39] = -15'd4389;
    value[40] = -15'd4386;
    value[41] = -15'd4383;
    value[42] = -15'd4380;
    value[43] = -15'd4377;
    value[44] = -15'd4374;
    value[45] = -15'd4371;
    value[46] = -15'd4368;
    value[47] = -15'd4365;
    value[48] = -15'd4363;
    value[49] = -15'd4360;
    value[50] = -15'd4357;
    value[51] = -15'd4354;
    value[52] = -15'd4351;
    value[53] = -15'd4348;
    value[54] = -15'd4345;
    value[55] = -15'd4342;
    value[56] = -15'd4339;
    value[57] = -15'd4336;
    value[58] = -15'd4333;
    value[59] = -15'd4330;
    value[60] = -15'd4327;
    value[61] = -15'd4324;
    value[62] = -15'd4321;
    value[63] = -15'd4318;
    value[64] = -15'd4315;
    value[65] = -15'd4312;
    value[66] = -15'd4309;
    value[67] = -15'd4306;
    value[68] = -15'd4303;
    value[69] = -15'd4300;
    value[70] = -15'd4297;
    value[71] = -15'd4294;
    value[72] = -15'd4291;
    value[73] = -15'd4288;
    value[74] = -15'd4285;
    value[75] = -15'd4282;
    value[76] = -15'd4279;
    value[77] = -15'd4276;
    value[78] = -15'd4273;
    value[79] = -15'd4270;
    value[80] = -15'd4267;
    value[81] = -15'd4264;
    value[82] = -15'd4261;
    value[83] = -15'd4258;
    value[84] = -15'd4255;
    value[85] = -15'd4252;
    value[86] = -15'd4249;
    value[87] = -15'd4246;
    value[88] = -15'd4243;
    value[89] = -15'd4240;
    value[90] = -15'd4237;
    value[91] = -15'd4234;
    value[92] = -15'd4231;
    value[93] = -15'd4228;
    value[94] = -15'd4225;
    value[95] = -15'd4222;
    value[96] = -15'd4218;
    value[97] = -15'd4215;
    value[98] = -15'd4212;
    value[99] = -15'd4209;
    value[100] = -15'd4206;
    value[101] = -15'd4203;
    value[102] = -15'd4200;
    value[103] = -15'd4197;
    value[104] = -15'd4194;
    value[105] = -15'd4191;
    value[106] = -15'd4188;
    value[107] = -15'd4184;
    value[108] = -15'd4181;
    value[109] = -15'd4178;
    value[110] = -15'd4175;
    value[111] = -15'd4172;
    value[112] = -15'd4169;
    value[113] = -15'd4166;
    value[114] = -15'd4163;
    value[115] = -15'd4160;
    value[116] = -15'd4156;
    value[117] = -15'd4153;
    value[118] = -15'd4150;
    value[119] = -15'd4147;
    value[120] = -15'd4144;
    value[121] = -15'd4141;
    value[122] = -15'd4138;
    value[123] = -15'd4134;
    value[124] = -15'd4131;
    value[125] = -15'd4128;
    value[126] = -15'd4125;
    value[127] = -15'd4122;
    value[128] = -15'd4119;
    value[129] = -15'd4115;
    value[130] = -15'd4112;
    value[131] = -15'd4109;
    value[132] = -15'd4106;
    value[133] = -15'd4103;
    value[134] = -15'd4100;
    value[135] = -15'd4096;
    value[136] = -15'd4093;
    value[137] = -15'd4090;
    value[138] = -15'd4087;
    value[139] = -15'd4084;
    value[140] = -15'd4080;
    value[141] = -15'd4077;
    value[142] = -15'd4074;
    value[143] = -15'd4071;
    value[144] = -15'd4067;
    value[145] = -15'd4064;
    value[146] = -15'd4061;
    value[147] = -15'd4058;
    value[148] = -15'd4055;
    value[149] = -15'd4051;
    value[150] = -15'd4048;
    value[151] = -15'd4045;
    value[152] = -15'd4042;
    value[153] = -15'd4038;
    value[154] = -15'd4035;
    value[155] = -15'd4032;
    value[156] = -15'd4029;
    value[157] = -15'd4025;
    value[158] = -15'd4022;
    value[159] = -15'd4019;
    value[160] = -15'd4016;
    value[161] = -15'd4012;
    value[162] = -15'd4009;
    value[163] = -15'd4006;
    value[164] = -15'd4003;
    value[165] = -15'd3999;
    value[166] = -15'd3996;
    value[167] = -15'd3993;
    value[168] = -15'd3989;
    value[169] = -15'd3986;
    value[170] = -15'd3983;
    value[171] = -15'd3979;
    value[172] = -15'd3976;
    value[173] = -15'd3973;
    value[174] = -15'd3970;
    value[175] = -15'd3966;
    value[176] = -15'd3963;
    value[177] = -15'd3960;
    value[178] = -15'd3956;
    value[179] = -15'd3953;
    value[180] = -15'd3950;
    value[181] = -15'd3946;
    value[182] = -15'd3943;
    value[183] = -15'd3940;
    value[184] = -15'd3936;
    value[185] = -15'd3933;
    value[186] = -15'd3930;
    value[187] = -15'd3926;
    value[188] = -15'd3923;
    value[189] = -15'd3919;
    value[190] = -15'd3916;
    value[191] = -15'd3913;
    value[192] = -15'd3909;
    value[193] = -15'd3906;
    value[194] = -15'd3903;
    value[195] = -15'd3899;
    value[196] = -15'd3896;
    value[197] = -15'd3892;
    value[198] = -15'd3889;
    value[199] = -15'd3886;
    value[200] = -15'd3882;
    value[201] = -15'd3879;
    value[202] = -15'd3876;
    value[203] = -15'd3872;
    value[204] = -15'd3869;
    value[205] = -15'd3865;
    value[206] = -15'd3862;
    value[207] = -15'd3858;
    value[208] = -15'd3855;
    value[209] = -15'd3852;
    value[210] = -15'd3848;
    value[211] = -15'd3845;
    value[212] = -15'd3841;
    value[213] = -15'd3838;
    value[214] = -15'd3834;
    value[215] = -15'd3831;
    value[216] = -15'd3828;
    value[217] = -15'd3824;
    value[218] = -15'd3821;
    value[219] = -15'd3817;
    value[220] = -15'd3814;
    value[221] = -15'd3810;
    value[222] = -15'd3807;
    value[223] = -15'd3803;
    value[224] = -15'd3800;
    value[225] = -15'd3796;
    value[226] = -15'd3793;
    value[227] = -15'd3789;
    value[228] = -15'd3786;
    value[229] = -15'd3782;
    value[230] = -15'd3779;
    value[231] = -15'd3775;
    value[232] = -15'd3772;
    value[233] = -15'd3768;
    value[234] = -15'd3765;
    value[235] = -15'd3761;
    value[236] = -15'd3758;
    value[237] = -15'd3754;
    value[238] = -15'd3751;
    value[239] = -15'd3747;
    value[240] = -15'd3744;
    value[241] = -15'd3740;
    value[242] = -15'd3737;
    value[243] = -15'd3733;
    value[244] = -15'd3730;
    value[245] = -15'd3726;
    value[246] = -15'd3723;
    value[247] = -15'd3719;
    value[248] = -15'd3716;
    value[249] = -15'd3712;
    value[250] = -15'd3708;
    value[251] = -15'd3705;
    value[252] = -15'd3701;
    value[253] = -15'd3698;
    value[254] = -15'd3694;
    value[255] = -15'd3691;
    value[256] = -15'd3687;
    value[257] = -15'd3683;
    value[258] = -15'd3680;
    value[259] = -15'd3676;
    value[260] = -15'd3673;
    value[261] = -15'd3669;
    value[262] = -15'd3665;
    value[263] = -15'd3662;
    value[264] = -15'd3658;
    value[265] = -15'd3655;
    value[266] = -15'd3651;
    value[267] = -15'd3647;
    value[268] = -15'd3644;
    value[269] = -15'd3640;
    value[270] = -15'd3637;
    value[271] = -15'd3633;
    value[272] = -15'd3629;
    value[273] = -15'd3626;
    value[274] = -15'd3622;
    value[275] = -15'd3618;
    value[276] = -15'd3615;
    value[277] = -15'd3611;
    value[278] = -15'd3607;
    value[279] = -15'd3604;
    value[280] = -15'd3600;
    value[281] = -15'd3596;
    value[282] = -15'd3593;
    value[283] = -15'd3589;
    value[284] = -15'd3585;
    value[285] = -15'd3582;
    value[286] = -15'd3578;
    value[287] = -15'd3574;
    value[288] = -15'd3571;
    value[289] = -15'd3567;
    value[290] = -15'd3563;
    value[291] = -15'd3560;
    value[292] = -15'd3556;
    value[293] = -15'd3552;
    value[294] = -15'd3548;
    value[295] = -15'd3545;
    value[296] = -15'd3541;
    value[297] = -15'd3537;
    value[298] = -15'd3534;
    value[299] = -15'd3530;
    value[300] = -15'd3526;
    value[301] = -15'd3522;
    value[302] = -15'd3519;
    value[303] = -15'd3515;
    value[304] = -15'd3511;
    value[305] = -15'd3507;
    value[306] = -15'd3504;
    value[307] = -15'd3500;
    value[308] = -15'd3496;
    value[309] = -15'd3492;
    value[310] = -15'd3489;
    value[311] = -15'd3485;
    value[312] = -15'd3481;
    value[313] = -15'd3477;
    value[314] = -15'd3474;
    value[315] = -15'd3470;
    value[316] = -15'd3466;
    value[317] = -15'd3462;
    value[318] = -15'd3458;
    value[319] = -15'd3455;
    value[320] = -15'd3451;
    value[321] = -15'd3447;
    value[322] = -15'd3443;
    value[323] = -15'd3439;
    value[324] = -15'd3436;
    value[325] = -15'd3432;
    value[326] = -15'd3428;
    value[327] = -15'd3424;
    value[328] = -15'd3420;
    value[329] = -15'd3417;
    value[330] = -15'd3413;
    value[331] = -15'd3409;
    value[332] = -15'd3405;
    value[333] = -15'd3401;
    value[334] = -15'd3397;
    value[335] = -15'd3393;
    value[336] = -15'd3390;
    value[337] = -15'd3386;
    value[338] = -15'd3382;
    value[339] = -15'd3378;
    value[340] = -15'd3374;
    value[341] = -15'd3370;
    value[342] = -15'd3366;
    value[343] = -15'd3363;
    value[344] = -15'd3359;
    value[345] = -15'd3355;
    value[346] = -15'd3351;
    value[347] = -15'd3347;
    value[348] = -15'd3343;
    value[349] = -15'd3339;
    value[350] = -15'd3335;
    value[351] = -15'd3331;
    value[352] = -15'd3327;
    value[353] = -15'd3324;
    value[354] = -15'd3320;
    value[355] = -15'd3316;
    value[356] = -15'd3312;
    value[357] = -15'd3308;
    value[358] = -15'd3304;
    value[359] = -15'd3300;
    value[360] = -15'd3296;
    value[361] = -15'd3292;
    value[362] = -15'd3288;
    value[363] = -15'd3284;
    value[364] = -15'd3280;
    value[365] = -15'd3276;
    value[366] = -15'd3272;
    value[367] = -15'd3268;
    value[368] = -15'd3264;
    value[369] = -15'd3260;
    value[370] = -15'd3257;
    value[371] = -15'd3253;
    value[372] = -15'd3249;
    value[373] = -15'd3245;
    value[374] = -15'd3241;
    value[375] = -15'd3237;
    value[376] = -15'd3233;
    value[377] = -15'd3229;
    value[378] = -15'd3225;
    value[379] = -15'd3221;
    value[380] = -15'd3217;
    value[381] = -15'd3213;
    value[382] = -15'd3209;
    value[383] = -15'd3205;
    value[384] = -15'd3201;
    value[385] = -15'd3197;
    value[386] = -15'd3192;
    value[387] = -15'd3188;
    value[388] = -15'd3184;
    value[389] = -15'd3180;
    value[390] = -15'd3176;
    value[391] = -15'd3172;
    value[392] = -15'd3168;
    value[393] = -15'd3164;
    value[394] = -15'd3160;
    value[395] = -15'd3156;
    value[396] = -15'd3152;
    value[397] = -15'd3148;
    value[398] = -15'd3144;
    value[399] = -15'd3140;
    value[400] = -15'd3136;
    value[401] = -15'd3132;
    value[402] = -15'd3128;
    value[403] = -15'd3123;
    value[404] = -15'd3119;
    value[405] = -15'd3115;
    value[406] = -15'd3111;
    value[407] = -15'd3107;
    value[408] = -15'd3103;
    value[409] = -15'd3099;
    value[410] = -15'd3095;
    value[411] = -15'd3091;
    value[412] = -15'd3086;
    value[413] = -15'd3082;
    value[414] = -15'd3078;
    value[415] = -15'd3074;
    value[416] = -15'd3070;
    value[417] = -15'd3066;
    value[418] = -15'd3062;
    value[419] = -15'd3058;
    value[420] = -15'd3053;
    value[421] = -15'd3049;
    value[422] = -15'd3045;
    value[423] = -15'd3041;
    value[424] = -15'd3037;
    value[425] = -15'd3033;
    value[426] = -15'd3028;
    value[427] = -15'd3024;
    value[428] = -15'd3020;
    value[429] = -15'd3016;
    value[430] = -15'd3012;
    value[431] = -15'd3008;
    value[432] = -15'd3003;
    value[433] = -15'd2999;
    value[434] = -15'd2995;
    value[435] = -15'd2991;
    value[436] = -15'd2987;
    value[437] = -15'd2982;
    value[438] = -15'd2978;
    value[439] = -15'd2974;
    value[440] = -15'd2970;
    value[441] = -15'd2965;
    value[442] = -15'd2961;
    value[443] = -15'd2957;
    value[444] = -15'd2953;
    value[445] = -15'd2949;
    value[446] = -15'd2944;
    value[447] = -15'd2940;
    value[448] = -15'd2936;
    value[449] = -15'd2932;
    value[450] = -15'd2927;
    value[451] = -15'd2923;
    value[452] = -15'd2919;
    value[453] = -15'd2914;
    value[454] = -15'd2910;
    value[455] = -15'd2906;
    value[456] = -15'd2902;
    value[457] = -15'd2897;
    value[458] = -15'd2893;
    value[459] = -15'd2889;
    value[460] = -15'd2885;
    value[461] = -15'd2880;
    value[462] = -15'd2876;
    value[463] = -15'd2872;
    value[464] = -15'd2867;
    value[465] = -15'd2863;
    value[466] = -15'd2859;
    value[467] = -15'd2854;
    value[468] = -15'd2850;
    value[469] = -15'd2846;
    value[470] = -15'd2841;
    value[471] = -15'd2837;
    value[472] = -15'd2833;
    value[473] = -15'd2828;
    value[474] = -15'd2824;
    value[475] = -15'd2820;
    value[476] = -15'd2815;
    value[477] = -15'd2811;
    value[478] = -15'd2807;
    value[479] = -15'd2802;
    value[480] = -15'd2798;
    value[481] = -15'd2794;
    value[482] = -15'd2789;
    value[483] = -15'd2785;
    value[484] = -15'd2780;
    value[485] = -15'd2776;
    value[486] = -15'd2772;
    value[487] = -15'd2767;
    value[488] = -15'd2763;
    value[489] = -15'd2759;
    value[490] = -15'd2754;
    value[491] = -15'd2750;
    value[492] = -15'd2745;
    value[493] = -15'd2741;
    value[494] = -15'd2737;
    value[495] = -15'd2732;
    value[496] = -15'd2728;
    value[497] = -15'd2723;
    value[498] = -15'd2719;
    value[499] = -15'd2714;
    value[500] = -15'd2710;
    value[501] = -15'd2706;
    value[502] = -15'd2701;
    value[503] = -15'd2697;
    value[504] = -15'd2692;
    value[505] = -15'd2688;
    value[506] = -15'd2683;
    value[507] = -15'd2679;
    value[508] = -15'd2674;
    value[509] = -15'd2670;
    value[510] = -15'd2665;
    value[511] = -15'd2661;
    value[512] = -15'd2657;
    value[513] = -15'd2652;
    value[514] = -15'd2648;
    value[515] = -15'd2643;
    value[516] = -15'd2639;
    value[517] = -15'd2634;
    value[518] = -15'd2630;
    value[519] = -15'd2625;
    value[520] = -15'd2621;
    value[521] = -15'd2616;
    value[522] = -15'd2612;
    value[523] = -15'd2607;
    value[524] = -15'd2603;
    value[525] = -15'd2598;
    value[526] = -15'd2593;
    value[527] = -15'd2589;
    value[528] = -15'd2584;
    value[529] = -15'd2580;
    value[530] = -15'd2575;
    value[531] = -15'd2571;
    value[532] = -15'd2566;
    value[533] = -15'd2562;
    value[534] = -15'd2557;
    value[535] = -15'd2553;
    value[536] = -15'd2548;
    value[537] = -15'd2544;
    value[538] = -15'd2539;
    value[539] = -15'd2534;
    value[540] = -15'd2530;
    value[541] = -15'd2525;
    value[542] = -15'd2521;
    value[543] = -15'd2516;
    value[544] = -15'd2511;
    value[545] = -15'd2507;
    value[546] = -15'd2502;
    value[547] = -15'd2498;
    value[548] = -15'd2493;
    value[549] = -15'd2489;
    value[550] = -15'd2484;
    value[551] = -15'd2479;
    value[552] = -15'd2475;
    value[553] = -15'd2470;
    value[554] = -15'd2465;
    value[555] = -15'd2461;
    value[556] = -15'd2456;
    value[557] = -15'd2452;
    value[558] = -15'd2447;
    value[559] = -15'd2442;
    value[560] = -15'd2438;
    value[561] = -15'd2433;
    value[562] = -15'd2428;
    value[563] = -15'd2424;
    value[564] = -15'd2419;
    value[565] = -15'd2414;
    value[566] = -15'd2410;
    value[567] = -15'd2405;
    value[568] = -15'd2400;
    value[569] = -15'd2396;
    value[570] = -15'd2391;
    value[571] = -15'd2386;
    value[572] = -15'd2382;
    value[573] = -15'd2377;
    value[574] = -15'd2372;
    value[575] = -15'd2368;
    value[576] = -15'd2363;
    value[577] = -15'd2358;
    value[578] = -15'd2354;
    value[579] = -15'd2349;
    value[580] = -15'd2344;
    value[581] = -15'd2339;
    value[582] = -15'd2335;
    value[583] = -15'd2330;
    value[584] = -15'd2325;
    value[585] = -15'd2321;
    value[586] = -15'd2316;
    value[587] = -15'd2311;
    value[588] = -15'd2306;
    value[589] = -15'd2302;
    value[590] = -15'd2297;
    value[591] = -15'd2292;
    value[592] = -15'd2287;
    value[593] = -15'd2283;
    value[594] = -15'd2278;
    value[595] = -15'd2273;
    value[596] = -15'd2268;
    value[597] = -15'd2264;
    value[598] = -15'd2259;
    value[599] = -15'd2254;
    value[600] = -15'd2249;
    value[601] = -15'd2244;
    value[602] = -15'd2240;
    value[603] = -15'd2235;
    value[604] = -15'd2230;
    value[605] = -15'd2225;
    value[606] = -15'd2221;
    value[607] = -15'd2216;
    value[608] = -15'd2211;
    value[609] = -15'd2206;
    value[610] = -15'd2201;
    value[611] = -15'd2197;
    value[612] = -15'd2192;
    value[613] = -15'd2187;
    value[614] = -15'd2182;
    value[615] = -15'd2177;
    value[616] = -15'd2172;
    value[617] = -15'd2168;
    value[618] = -15'd2163;
    value[619] = -15'd2158;
    value[620] = -15'd2153;
    value[621] = -15'd2148;
    value[622] = -15'd2143;
    value[623] = -15'd2139;
    value[624] = -15'd2134;
    value[625] = -15'd2129;
    value[626] = -15'd2124;
    value[627] = -15'd2119;
    value[628] = -15'd2114;
    value[629] = -15'd2109;
    value[630] = -15'd2105;
    value[631] = -15'd2100;
    value[632] = -15'd2095;
    value[633] = -15'd2090;
    value[634] = -15'd2085;
    value[635] = -15'd2080;
    value[636] = -15'd2075;
    value[637] = -15'd2070;
    value[638] = -15'd2065;
    value[639] = -15'd2061;
    value[640] = -15'd2056;
    value[641] = -15'd2051;
    value[642] = -15'd2046;
    value[643] = -15'd2041;
    value[644] = -15'd2036;
    value[645] = -15'd2031;
    value[646] = -15'd2026;
    value[647] = -15'd2021;
    value[648] = -15'd2016;
    value[649] = -15'd2011;
    value[650] = -15'd2006;
    value[651] = -15'd2001;
    value[652] = -15'd1997;
    value[653] = -15'd1992;
    value[654] = -15'd1987;
    value[655] = -15'd1982;
    value[656] = -15'd1977;
    value[657] = -15'd1972;
    value[658] = -15'd1967;
    value[659] = -15'd1962;
    value[660] = -15'd1957;
    value[661] = -15'd1952;
    value[662] = -15'd1947;
    value[663] = -15'd1942;
    value[664] = -15'd1937;
    value[665] = -15'd1932;
    value[666] = -15'd1927;
    value[667] = -15'd1922;
    value[668] = -15'd1917;
    value[669] = -15'd1912;
    value[670] = -15'd1907;
    value[671] = -15'd1902;
    value[672] = -15'd1897;
    value[673] = -15'd1892;
    value[674] = -15'd1887;
    value[675] = -15'd1882;
    value[676] = -15'd1877;
    value[677] = -15'd1872;
    value[678] = -15'd1867;
    value[679] = -15'd1862;
    value[680] = -15'd1857;
    value[681] = -15'd1852;
    value[682] = -15'd1847;
    value[683] = -15'd1842;
    value[684] = -15'd1837;
    value[685] = -15'd1832;
    value[686] = -15'd1827;
    value[687] = -15'd1822;
    value[688] = -15'd1817;
    value[689] = -15'd1812;
    value[690] = -15'd1806;
    value[691] = -15'd1801;
    value[692] = -15'd1796;
    value[693] = -15'd1791;
    value[694] = -15'd1786;
    value[695] = -15'd1781;
    value[696] = -15'd1776;
    value[697] = -15'd1771;
    value[698] = -15'd1766;
    value[699] = -15'd1761;
    value[700] = -15'd1756;
    value[701] = -15'd1751;
    value[702] = -15'd1746;
    value[703] = -15'd1740;
    value[704] = -15'd1735;
    value[705] = -15'd1730;
    value[706] = -15'd1725;
    value[707] = -15'd1720;
    value[708] = -15'd1715;
    value[709] = -15'd1710;
    value[710] = -15'd1705;
    value[711] = -15'd1700;
    value[712] = -15'd1695;
    value[713] = -15'd1689;
    value[714] = -15'd1684;
    value[715] = -15'd1679;
    value[716] = -15'd1674;
    value[717] = -15'd1669;
    value[718] = -15'd1664;
    value[719] = -15'd1659;
    value[720] = -15'd1653;
    value[721] = -15'd1648;
    value[722] = -15'd1643;
    value[723] = -15'd1638;
    value[724] = -15'd1633;
    value[725] = -15'd1628;
    value[726] = -15'd1623;
    value[727] = -15'd1617;
    value[728] = -15'd1612;
    value[729] = -15'd1607;
    value[730] = -15'd1602;
    value[731] = -15'd1597;
    value[732] = -15'd1592;
    value[733] = -15'd1586;
    value[734] = -15'd1581;
    value[735] = -15'd1576;
    value[736] = -15'd1571;
    value[737] = -15'd1566;
    value[738] = -15'd1560;
    value[739] = -15'd1555;
    value[740] = -15'd1550;
    value[741] = -15'd1545;
    value[742] = -15'd1540;
    value[743] = -15'd1535;
    value[744] = -15'd1529;
    value[745] = -15'd1524;
    value[746] = -15'd1519;
    value[747] = -15'd1514;
    value[748] = -15'd1508;
    value[749] = -15'd1503;
    value[750] = -15'd1498;
    value[751] = -15'd1493;
    value[752] = -15'd1488;
    value[753] = -15'd1482;
    value[754] = -15'd1477;
    value[755] = -15'd1472;
    value[756] = -15'd1467;
    value[757] = -15'd1461;
    value[758] = -15'd1456;
    value[759] = -15'd1451;
    value[760] = -15'd1446;
    value[761] = -15'd1440;
    value[762] = -15'd1435;
    value[763] = -15'd1430;
    value[764] = -15'd1425;
    value[765] = -15'd1419;
    value[766] = -15'd1414;
    value[767] = -15'd1409;
    value[768] = -15'd1404;
    value[769] = -15'd1398;
    value[770] = -15'd1393;
    value[771] = -15'd1388;
    value[772] = -15'd1383;
    value[773] = -15'd1377;
    value[774] = -15'd1372;
    value[775] = -15'd1367;
    value[776] = -15'd1361;
    value[777] = -15'd1356;
    value[778] = -15'd1351;
    value[779] = -15'd1346;
    value[780] = -15'd1340;
    value[781] = -15'd1335;
    value[782] = -15'd1330;
    value[783] = -15'd1324;
    value[784] = -15'd1319;
    value[785] = -15'd1314;
    value[786] = -15'd1308;
    value[787] = -15'd1303;
    value[788] = -15'd1298;
    value[789] = -15'd1293;
    value[790] = -15'd1287;
    value[791] = -15'd1282;
    value[792] = -15'd1277;
    value[793] = -15'd1271;
    value[794] = -15'd1266;
    value[795] = -15'd1261;
    value[796] = -15'd1255;
    value[797] = -15'd1250;
    value[798] = -15'd1245;
    value[799] = -15'd1239;
    value[800] = -15'd1234;
    value[801] = -15'd1229;
    value[802] = -15'd1223;
    value[803] = -15'd1218;
    value[804] = -15'd1213;
    value[805] = -15'd1207;
    value[806] = -15'd1202;
    value[807] = -15'd1196;
    value[808] = -15'd1191;
    value[809] = -15'd1186;
    value[810] = -15'd1180;
    value[811] = -15'd1175;
    value[812] = -15'd1170;
    value[813] = -15'd1164;
    value[814] = -15'd1159;
    value[815] = -15'd1154;
    value[816] = -15'd1148;
    value[817] = -15'd1143;
    value[818] = -15'd1137;
    value[819] = -15'd1132;
    value[820] = -15'd1127;
    value[821] = -15'd1121;
    value[822] = -15'd1116;
    value[823] = -15'd1111;
    value[824] = -15'd1105;
    value[825] = -15'd1100;
    value[826] = -15'd1094;
    value[827] = -15'd1089;
    value[828] = -15'd1084;
    value[829] = -15'd1078;
    value[830] = -15'd1073;
    value[831] = -15'd1067;
    value[832] = -15'd1062;
    value[833] = -15'd1057;
    value[834] = -15'd1051;
    value[835] = -15'd1046;
    value[836] = -15'd1040;
    value[837] = -15'd1035;
    value[838] = -15'd1029;
    value[839] = -15'd1024;
    value[840] = -15'd1019;
    value[841] = -15'd1013;
    value[842] = -15'd1008;
    value[843] = -15'd1002;
    value[844] = -15'd997;
    value[845] = -15'd992;
    value[846] = -15'd986;
    value[847] = -15'd981;
    value[848] = -15'd975;
    value[849] = -15'd970;
    value[850] = -15'd964;
    value[851] = -15'd959;
    value[852] = -15'd953;
    value[853] = -15'd948;
    value[854] = -15'd943;
    value[855] = -15'd937;
    value[856] = -15'd932;
    value[857] = -15'd926;
    value[858] = -15'd921;
    value[859] = -15'd915;
    value[860] = -15'd910;
    value[861] = -15'd904;
    value[862] = -15'd899;
    value[863] = -15'd894;
    value[864] = -15'd888;
    value[865] = -15'd883;
    value[866] = -15'd877;
    value[867] = -15'd872;
    value[868] = -15'd866;
    value[869] = -15'd861;
    value[870] = -15'd855;
    value[871] = -15'd850;
    value[872] = -15'd844;
    value[873] = -15'd839;
    value[874] = -15'd833;
    value[875] = -15'd828;
    value[876] = -15'd822;
    value[877] = -15'd817;
    value[878] = -15'd811;
    value[879] = -15'd806;
    value[880] = -15'd800;
    value[881] = -15'd795;
    value[882] = -15'd789;
    value[883] = -15'd784;
    value[884] = -15'd779;
    value[885] = -15'd773;
    value[886] = -15'd768;
    value[887] = -15'd762;
    value[888] = -15'd757;
    value[889] = -15'd751;
    value[890] = -15'd746;
    value[891] = -15'd740;
    value[892] = -15'd735;
    value[893] = -15'd729;
    value[894] = -15'd724;
    value[895] = -15'd718;
    value[896] = -15'd713;
    value[897] = -15'd707;
    value[898] = -15'd701;
    value[899] = -15'd696;
    value[900] = -15'd690;
    value[901] = -15'd685;
    value[902] = -15'd679;
    value[903] = -15'd674;
    value[904] = -15'd668;
    value[905] = -15'd663;
    value[906] = -15'd657;
    value[907] = -15'd652;
    value[908] = -15'd646;
    value[909] = -15'd641;
    value[910] = -15'd635;
    value[911] = -15'd630;
    value[912] = -15'd624;
    value[913] = -15'd619;
    value[914] = -15'd613;
    value[915] = -15'd608;
    value[916] = -15'd602;
    value[917] = -15'd597;
    value[918] = -15'd591;
    value[919] = -15'd585;
    value[920] = -15'd580;
    value[921] = -15'd574;
    value[922] = -15'd569;
    value[923] = -15'd563;
    value[924] = -15'd558;
    value[925] = -15'd552;
    value[926] = -15'd547;
    value[927] = -15'd541;
    value[928] = -15'd536;
    value[929] = -15'd530;
    value[930] = -15'd524;
    value[931] = -15'd519;
    value[932] = -15'd513;
    value[933] = -15'd508;
    value[934] = -15'd502;
    value[935] = -15'd497;
    value[936] = -15'd491;
    value[937] = -15'd486;
    value[938] = -15'd480;
    value[939] = -15'd475;
    value[940] = -15'd469;
    value[941] = -15'd463;
    value[942] = -15'd458;
    value[943] = -15'd452;
    value[944] = -15'd447;
    value[945] = -15'd441;
    value[946] = -15'd436;
    value[947] = -15'd430;
    value[948] = -15'd424;
    value[949] = -15'd419;
    value[950] = -15'd413;
    value[951] = -15'd408;
    value[952] = -15'd402;
    value[953] = -15'd397;
    value[954] = -15'd391;
    value[955] = -15'd385;
    value[956] = -15'd380;
    value[957] = -15'd374;
    value[958] = -15'd369;
    value[959] = -15'd363;
    value[960] = -15'd358;
    value[961] = -15'd352;
    value[962] = -15'd346;
    value[963] = -15'd341;
    value[964] = -15'd335;
    value[965] = -15'd330;
    value[966] = -15'd324;
    value[967] = -15'd319;
    value[968] = -15'd313;
    value[969] = -15'd307;
    value[970] = -15'd302;
    value[971] = -15'd296;
    value[972] = -15'd291;
    value[973] = -15'd285;
    value[974] = -15'd280;
    value[975] = -15'd274;
    value[976] = -15'd268;
    value[977] = -15'd263;
    value[978] = -15'd257;
    value[979] = -15'd252;
    value[980] = -15'd246;
    value[981] = -15'd240;
    value[982] = -15'd235;
    value[983] = -15'd229;
    value[984] = -15'd224;
    value[985] = -15'd218;
    value[986] = -15'd213;
    value[987] = -15'd207;
    value[988] = -15'd201;
    value[989] = -15'd196;
    value[990] = -15'd190;
    value[991] = -15'd185;
    value[992] = -15'd179;
    value[993] = -15'd173;
    value[994] = -15'd168;
    value[995] = -15'd162;
    value[996] = -15'd157;
    value[997] = -15'd151;
    value[998] = -15'd145;
    value[999] = -15'd140;
    value[1000] = -15'd134;
    value[1001] = -15'd129;
    value[1002] = -15'd123;
    value[1003] = -15'd117;
    value[1004] = -15'd112;
    value[1005] = -15'd106;
    value[1006] = -15'd101;
    value[1007] = -15'd95;
    value[1008] = -15'd90;
    value[1009] = -15'd84;
    value[1010] = -15'd78;
    value[1011] = -15'd73;
    value[1012] = -15'd67;
    value[1013] = -15'd62;
    value[1014] = -15'd56;
    value[1015] = -15'd50;
    value[1016] = -15'd45;
    value[1017] = -15'd39;
    value[1018] = -15'd34;
    value[1019] = -15'd28;
    value[1020] = -15'd22;
    value[1021] = -15'd17;
    value[1022] = -15'd11;
    value[1023] = -15'd6;
    value[1024] = 15'd0;
    value[1025] = 15'd6;
    value[1026] = 15'd11;
    value[1027] = 15'd17;
    value[1028] = 15'd22;
    value[1029] = 15'd28;
    value[1030] = 15'd34;
    value[1031] = 15'd39;
    value[1032] = 15'd45;
    value[1033] = 15'd50;
    value[1034] = 15'd56;
    value[1035] = 15'd62;
    value[1036] = 15'd67;
    value[1037] = 15'd73;
    value[1038] = 15'd78;
    value[1039] = 15'd84;
    value[1040] = 15'd90;
    value[1041] = 15'd95;
    value[1042] = 15'd101;
    value[1043] = 15'd106;
    value[1044] = 15'd112;
    value[1045] = 15'd117;
    value[1046] = 15'd123;
    value[1047] = 15'd129;
    value[1048] = 15'd134;
    value[1049] = 15'd140;
    value[1050] = 15'd145;
    value[1051] = 15'd151;
    value[1052] = 15'd157;
    value[1053] = 15'd162;
    value[1054] = 15'd168;
    value[1055] = 15'd173;
    value[1056] = 15'd179;
    value[1057] = 15'd185;
    value[1058] = 15'd190;
    value[1059] = 15'd196;
    value[1060] = 15'd201;
    value[1061] = 15'd207;
    value[1062] = 15'd213;
    value[1063] = 15'd218;
    value[1064] = 15'd224;
    value[1065] = 15'd229;
    value[1066] = 15'd235;
    value[1067] = 15'd240;
    value[1068] = 15'd246;
    value[1069] = 15'd252;
    value[1070] = 15'd257;
    value[1071] = 15'd263;
    value[1072] = 15'd268;
    value[1073] = 15'd274;
    value[1074] = 15'd280;
    value[1075] = 15'd285;
    value[1076] = 15'd291;
    value[1077] = 15'd296;
    value[1078] = 15'd302;
    value[1079] = 15'd307;
    value[1080] = 15'd313;
    value[1081] = 15'd319;
    value[1082] = 15'd324;
    value[1083] = 15'd330;
    value[1084] = 15'd335;
    value[1085] = 15'd341;
    value[1086] = 15'd346;
    value[1087] = 15'd352;
    value[1088] = 15'd358;
    value[1089] = 15'd363;
    value[1090] = 15'd369;
    value[1091] = 15'd374;
    value[1092] = 15'd380;
    value[1093] = 15'd385;
    value[1094] = 15'd391;
    value[1095] = 15'd397;
    value[1096] = 15'd402;
    value[1097] = 15'd408;
    value[1098] = 15'd413;
    value[1099] = 15'd419;
    value[1100] = 15'd424;
    value[1101] = 15'd430;
    value[1102] = 15'd436;
    value[1103] = 15'd441;
    value[1104] = 15'd447;
    value[1105] = 15'd452;
    value[1106] = 15'd458;
    value[1107] = 15'd463;
    value[1108] = 15'd469;
    value[1109] = 15'd475;
    value[1110] = 15'd480;
    value[1111] = 15'd486;
    value[1112] = 15'd491;
    value[1113] = 15'd497;
    value[1114] = 15'd502;
    value[1115] = 15'd508;
    value[1116] = 15'd513;
    value[1117] = 15'd519;
    value[1118] = 15'd524;
    value[1119] = 15'd530;
    value[1120] = 15'd536;
    value[1121] = 15'd541;
    value[1122] = 15'd547;
    value[1123] = 15'd552;
    value[1124] = 15'd558;
    value[1125] = 15'd563;
    value[1126] = 15'd569;
    value[1127] = 15'd574;
    value[1128] = 15'd580;
    value[1129] = 15'd585;
    value[1130] = 15'd591;
    value[1131] = 15'd597;
    value[1132] = 15'd602;
    value[1133] = 15'd608;
    value[1134] = 15'd613;
    value[1135] = 15'd619;
    value[1136] = 15'd624;
    value[1137] = 15'd630;
    value[1138] = 15'd635;
    value[1139] = 15'd641;
    value[1140] = 15'd646;
    value[1141] = 15'd652;
    value[1142] = 15'd657;
    value[1143] = 15'd663;
    value[1144] = 15'd668;
    value[1145] = 15'd674;
    value[1146] = 15'd679;
    value[1147] = 15'd685;
    value[1148] = 15'd690;
    value[1149] = 15'd696;
    value[1150] = 15'd701;
    value[1151] = 15'd707;
    value[1152] = 15'd713;
    value[1153] = 15'd718;
    value[1154] = 15'd724;
    value[1155] = 15'd729;
    value[1156] = 15'd735;
    value[1157] = 15'd740;
    value[1158] = 15'd746;
    value[1159] = 15'd751;
    value[1160] = 15'd757;
    value[1161] = 15'd762;
    value[1162] = 15'd768;
    value[1163] = 15'd773;
    value[1164] = 15'd779;
    value[1165] = 15'd784;
    value[1166] = 15'd789;
    value[1167] = 15'd795;
    value[1168] = 15'd800;
    value[1169] = 15'd806;
    value[1170] = 15'd811;
    value[1171] = 15'd817;
    value[1172] = 15'd822;
    value[1173] = 15'd828;
    value[1174] = 15'd833;
    value[1175] = 15'd839;
    value[1176] = 15'd844;
    value[1177] = 15'd850;
    value[1178] = 15'd855;
    value[1179] = 15'd861;
    value[1180] = 15'd866;
    value[1181] = 15'd872;
    value[1182] = 15'd877;
    value[1183] = 15'd883;
    value[1184] = 15'd888;
    value[1185] = 15'd894;
    value[1186] = 15'd899;
    value[1187] = 15'd904;
    value[1188] = 15'd910;
    value[1189] = 15'd915;
    value[1190] = 15'd921;
    value[1191] = 15'd926;
    value[1192] = 15'd932;
    value[1193] = 15'd937;
    value[1194] = 15'd943;
    value[1195] = 15'd948;
    value[1196] = 15'd953;
    value[1197] = 15'd959;
    value[1198] = 15'd964;
    value[1199] = 15'd970;
    value[1200] = 15'd975;
    value[1201] = 15'd981;
    value[1202] = 15'd986;
    value[1203] = 15'd992;
    value[1204] = 15'd997;
    value[1205] = 15'd1002;
    value[1206] = 15'd1008;
    value[1207] = 15'd1013;
    value[1208] = 15'd1019;
    value[1209] = 15'd1024;
    value[1210] = 15'd1029;
    value[1211] = 15'd1035;
    value[1212] = 15'd1040;
    value[1213] = 15'd1046;
    value[1214] = 15'd1051;
    value[1215] = 15'd1057;
    value[1216] = 15'd1062;
    value[1217] = 15'd1067;
    value[1218] = 15'd1073;
    value[1219] = 15'd1078;
    value[1220] = 15'd1084;
    value[1221] = 15'd1089;
    value[1222] = 15'd1094;
    value[1223] = 15'd1100;
    value[1224] = 15'd1105;
    value[1225] = 15'd1111;
    value[1226] = 15'd1116;
    value[1227] = 15'd1121;
    value[1228] = 15'd1127;
    value[1229] = 15'd1132;
    value[1230] = 15'd1137;
    value[1231] = 15'd1143;
    value[1232] = 15'd1148;
    value[1233] = 15'd1154;
    value[1234] = 15'd1159;
    value[1235] = 15'd1164;
    value[1236] = 15'd1170;
    value[1237] = 15'd1175;
    value[1238] = 15'd1180;
    value[1239] = 15'd1186;
    value[1240] = 15'd1191;
    value[1241] = 15'd1196;
    value[1242] = 15'd1202;
    value[1243] = 15'd1207;
    value[1244] = 15'd1213;
    value[1245] = 15'd1218;
    value[1246] = 15'd1223;
    value[1247] = 15'd1229;
    value[1248] = 15'd1234;
    value[1249] = 15'd1239;
    value[1250] = 15'd1245;
    value[1251] = 15'd1250;
    value[1252] = 15'd1255;
    value[1253] = 15'd1261;
    value[1254] = 15'd1266;
    value[1255] = 15'd1271;
    value[1256] = 15'd1277;
    value[1257] = 15'd1282;
    value[1258] = 15'd1287;
    value[1259] = 15'd1293;
    value[1260] = 15'd1298;
    value[1261] = 15'd1303;
    value[1262] = 15'd1308;
    value[1263] = 15'd1314;
    value[1264] = 15'd1319;
    value[1265] = 15'd1324;
    value[1266] = 15'd1330;
    value[1267] = 15'd1335;
    value[1268] = 15'd1340;
    value[1269] = 15'd1346;
    value[1270] = 15'd1351;
    value[1271] = 15'd1356;
    value[1272] = 15'd1361;
    value[1273] = 15'd1367;
    value[1274] = 15'd1372;
    value[1275] = 15'd1377;
    value[1276] = 15'd1383;
    value[1277] = 15'd1388;
    value[1278] = 15'd1393;
    value[1279] = 15'd1398;
    value[1280] = 15'd1404;
    value[1281] = 15'd1409;
    value[1282] = 15'd1414;
    value[1283] = 15'd1419;
    value[1284] = 15'd1425;
    value[1285] = 15'd1430;
    value[1286] = 15'd1435;
    value[1287] = 15'd1440;
    value[1288] = 15'd1446;
    value[1289] = 15'd1451;
    value[1290] = 15'd1456;
    value[1291] = 15'd1461;
    value[1292] = 15'd1467;
    value[1293] = 15'd1472;
    value[1294] = 15'd1477;
    value[1295] = 15'd1482;
    value[1296] = 15'd1488;
    value[1297] = 15'd1493;
    value[1298] = 15'd1498;
    value[1299] = 15'd1503;
    value[1300] = 15'd1508;
    value[1301] = 15'd1514;
    value[1302] = 15'd1519;
    value[1303] = 15'd1524;
    value[1304] = 15'd1529;
    value[1305] = 15'd1535;
    value[1306] = 15'd1540;
    value[1307] = 15'd1545;
    value[1308] = 15'd1550;
    value[1309] = 15'd1555;
    value[1310] = 15'd1560;
    value[1311] = 15'd1566;
    value[1312] = 15'd1571;
    value[1313] = 15'd1576;
    value[1314] = 15'd1581;
    value[1315] = 15'd1586;
    value[1316] = 15'd1592;
    value[1317] = 15'd1597;
    value[1318] = 15'd1602;
    value[1319] = 15'd1607;
    value[1320] = 15'd1612;
    value[1321] = 15'd1617;
    value[1322] = 15'd1623;
    value[1323] = 15'd1628;
    value[1324] = 15'd1633;
    value[1325] = 15'd1638;
    value[1326] = 15'd1643;
    value[1327] = 15'd1648;
    value[1328] = 15'd1653;
    value[1329] = 15'd1659;
    value[1330] = 15'd1664;
    value[1331] = 15'd1669;
    value[1332] = 15'd1674;
    value[1333] = 15'd1679;
    value[1334] = 15'd1684;
    value[1335] = 15'd1689;
    value[1336] = 15'd1695;
    value[1337] = 15'd1700;
    value[1338] = 15'd1705;
    value[1339] = 15'd1710;
    value[1340] = 15'd1715;
    value[1341] = 15'd1720;
    value[1342] = 15'd1725;
    value[1343] = 15'd1730;
    value[1344] = 15'd1735;
    value[1345] = 15'd1740;
    value[1346] = 15'd1746;
    value[1347] = 15'd1751;
    value[1348] = 15'd1756;
    value[1349] = 15'd1761;
    value[1350] = 15'd1766;
    value[1351] = 15'd1771;
    value[1352] = 15'd1776;
    value[1353] = 15'd1781;
    value[1354] = 15'd1786;
    value[1355] = 15'd1791;
    value[1356] = 15'd1796;
    value[1357] = 15'd1801;
    value[1358] = 15'd1806;
    value[1359] = 15'd1812;
    value[1360] = 15'd1817;
    value[1361] = 15'd1822;
    value[1362] = 15'd1827;
    value[1363] = 15'd1832;
    value[1364] = 15'd1837;
    value[1365] = 15'd1842;
    value[1366] = 15'd1847;
    value[1367] = 15'd1852;
    value[1368] = 15'd1857;
    value[1369] = 15'd1862;
    value[1370] = 15'd1867;
    value[1371] = 15'd1872;
    value[1372] = 15'd1877;
    value[1373] = 15'd1882;
    value[1374] = 15'd1887;
    value[1375] = 15'd1892;
    value[1376] = 15'd1897;
    value[1377] = 15'd1902;
    value[1378] = 15'd1907;
    value[1379] = 15'd1912;
    value[1380] = 15'd1917;
    value[1381] = 15'd1922;
    value[1382] = 15'd1927;
    value[1383] = 15'd1932;
    value[1384] = 15'd1937;
    value[1385] = 15'd1942;
    value[1386] = 15'd1947;
    value[1387] = 15'd1952;
    value[1388] = 15'd1957;
    value[1389] = 15'd1962;
    value[1390] = 15'd1967;
    value[1391] = 15'd1972;
    value[1392] = 15'd1977;
    value[1393] = 15'd1982;
    value[1394] = 15'd1987;
    value[1395] = 15'd1992;
    value[1396] = 15'd1997;
    value[1397] = 15'd2001;
    value[1398] = 15'd2006;
    value[1399] = 15'd2011;
    value[1400] = 15'd2016;
    value[1401] = 15'd2021;
    value[1402] = 15'd2026;
    value[1403] = 15'd2031;
    value[1404] = 15'd2036;
    value[1405] = 15'd2041;
    value[1406] = 15'd2046;
    value[1407] = 15'd2051;
    value[1408] = 15'd2056;
    value[1409] = 15'd2061;
    value[1410] = 15'd2065;
    value[1411] = 15'd2070;
    value[1412] = 15'd2075;
    value[1413] = 15'd2080;
    value[1414] = 15'd2085;
    value[1415] = 15'd2090;
    value[1416] = 15'd2095;
    value[1417] = 15'd2100;
    value[1418] = 15'd2105;
    value[1419] = 15'd2109;
    value[1420] = 15'd2114;
    value[1421] = 15'd2119;
    value[1422] = 15'd2124;
    value[1423] = 15'd2129;
    value[1424] = 15'd2134;
    value[1425] = 15'd2139;
    value[1426] = 15'd2143;
    value[1427] = 15'd2148;
    value[1428] = 15'd2153;
    value[1429] = 15'd2158;
    value[1430] = 15'd2163;
    value[1431] = 15'd2168;
    value[1432] = 15'd2172;
    value[1433] = 15'd2177;
    value[1434] = 15'd2182;
    value[1435] = 15'd2187;
    value[1436] = 15'd2192;
    value[1437] = 15'd2197;
    value[1438] = 15'd2201;
    value[1439] = 15'd2206;
    value[1440] = 15'd2211;
    value[1441] = 15'd2216;
    value[1442] = 15'd2221;
    value[1443] = 15'd2225;
    value[1444] = 15'd2230;
    value[1445] = 15'd2235;
    value[1446] = 15'd2240;
    value[1447] = 15'd2244;
    value[1448] = 15'd2249;
    value[1449] = 15'd2254;
    value[1450] = 15'd2259;
    value[1451] = 15'd2264;
    value[1452] = 15'd2268;
    value[1453] = 15'd2273;
    value[1454] = 15'd2278;
    value[1455] = 15'd2283;
    value[1456] = 15'd2287;
    value[1457] = 15'd2292;
    value[1458] = 15'd2297;
    value[1459] = 15'd2302;
    value[1460] = 15'd2306;
    value[1461] = 15'd2311;
    value[1462] = 15'd2316;
    value[1463] = 15'd2321;
    value[1464] = 15'd2325;
    value[1465] = 15'd2330;
    value[1466] = 15'd2335;
    value[1467] = 15'd2339;
    value[1468] = 15'd2344;
    value[1469] = 15'd2349;
    value[1470] = 15'd2354;
    value[1471] = 15'd2358;
    value[1472] = 15'd2363;
    value[1473] = 15'd2368;
    value[1474] = 15'd2372;
    value[1475] = 15'd2377;
    value[1476] = 15'd2382;
    value[1477] = 15'd2386;
    value[1478] = 15'd2391;
    value[1479] = 15'd2396;
    value[1480] = 15'd2400;
    value[1481] = 15'd2405;
    value[1482] = 15'd2410;
    value[1483] = 15'd2414;
    value[1484] = 15'd2419;
    value[1485] = 15'd2424;
    value[1486] = 15'd2428;
    value[1487] = 15'd2433;
    value[1488] = 15'd2438;
    value[1489] = 15'd2442;
    value[1490] = 15'd2447;
    value[1491] = 15'd2452;
    value[1492] = 15'd2456;
    value[1493] = 15'd2461;
    value[1494] = 15'd2465;
    value[1495] = 15'd2470;
    value[1496] = 15'd2475;
    value[1497] = 15'd2479;
    value[1498] = 15'd2484;
    value[1499] = 15'd2489;
    value[1500] = 15'd2493;
    value[1501] = 15'd2498;
    value[1502] = 15'd2502;
    value[1503] = 15'd2507;
    value[1504] = 15'd2511;
    value[1505] = 15'd2516;
    value[1506] = 15'd2521;
    value[1507] = 15'd2525;
    value[1508] = 15'd2530;
    value[1509] = 15'd2534;
    value[1510] = 15'd2539;
    value[1511] = 15'd2544;
    value[1512] = 15'd2548;
    value[1513] = 15'd2553;
    value[1514] = 15'd2557;
    value[1515] = 15'd2562;
    value[1516] = 15'd2566;
    value[1517] = 15'd2571;
    value[1518] = 15'd2575;
    value[1519] = 15'd2580;
    value[1520] = 15'd2584;
    value[1521] = 15'd2589;
    value[1522] = 15'd2593;
    value[1523] = 15'd2598;
    value[1524] = 15'd2603;
    value[1525] = 15'd2607;
    value[1526] = 15'd2612;
    value[1527] = 15'd2616;
    value[1528] = 15'd2621;
    value[1529] = 15'd2625;
    value[1530] = 15'd2630;
    value[1531] = 15'd2634;
    value[1532] = 15'd2639;
    value[1533] = 15'd2643;
    value[1534] = 15'd2648;
    value[1535] = 15'd2652;
    value[1536] = 15'd2657;
    value[1537] = 15'd2661;
    value[1538] = 15'd2665;
    value[1539] = 15'd2670;
    value[1540] = 15'd2674;
    value[1541] = 15'd2679;
    value[1542] = 15'd2683;
    value[1543] = 15'd2688;
    value[1544] = 15'd2692;
    value[1545] = 15'd2697;
    value[1546] = 15'd2701;
    value[1547] = 15'd2706;
    value[1548] = 15'd2710;
    value[1549] = 15'd2714;
    value[1550] = 15'd2719;
    value[1551] = 15'd2723;
    value[1552] = 15'd2728;
    value[1553] = 15'd2732;
    value[1554] = 15'd2737;
    value[1555] = 15'd2741;
    value[1556] = 15'd2745;
    value[1557] = 15'd2750;
    value[1558] = 15'd2754;
    value[1559] = 15'd2759;
    value[1560] = 15'd2763;
    value[1561] = 15'd2767;
    value[1562] = 15'd2772;
    value[1563] = 15'd2776;
    value[1564] = 15'd2780;
    value[1565] = 15'd2785;
    value[1566] = 15'd2789;
    value[1567] = 15'd2794;
    value[1568] = 15'd2798;
    value[1569] = 15'd2802;
    value[1570] = 15'd2807;
    value[1571] = 15'd2811;
    value[1572] = 15'd2815;
    value[1573] = 15'd2820;
    value[1574] = 15'd2824;
    value[1575] = 15'd2828;
    value[1576] = 15'd2833;
    value[1577] = 15'd2837;
    value[1578] = 15'd2841;
    value[1579] = 15'd2846;
    value[1580] = 15'd2850;
    value[1581] = 15'd2854;
    value[1582] = 15'd2859;
    value[1583] = 15'd2863;
    value[1584] = 15'd2867;
    value[1585] = 15'd2872;
    value[1586] = 15'd2876;
    value[1587] = 15'd2880;
    value[1588] = 15'd2885;
    value[1589] = 15'd2889;
    value[1590] = 15'd2893;
    value[1591] = 15'd2897;
    value[1592] = 15'd2902;
    value[1593] = 15'd2906;
    value[1594] = 15'd2910;
    value[1595] = 15'd2914;
    value[1596] = 15'd2919;
    value[1597] = 15'd2923;
    value[1598] = 15'd2927;
    value[1599] = 15'd2932;
    value[1600] = 15'd2936;
    value[1601] = 15'd2940;
    value[1602] = 15'd2944;
    value[1603] = 15'd2949;
    value[1604] = 15'd2953;
    value[1605] = 15'd2957;
    value[1606] = 15'd2961;
    value[1607] = 15'd2965;
    value[1608] = 15'd2970;
    value[1609] = 15'd2974;
    value[1610] = 15'd2978;
    value[1611] = 15'd2982;
    value[1612] = 15'd2987;
    value[1613] = 15'd2991;
    value[1614] = 15'd2995;
    value[1615] = 15'd2999;
    value[1616] = 15'd3003;
    value[1617] = 15'd3008;
    value[1618] = 15'd3012;
    value[1619] = 15'd3016;
    value[1620] = 15'd3020;
    value[1621] = 15'd3024;
    value[1622] = 15'd3028;
    value[1623] = 15'd3033;
    value[1624] = 15'd3037;
    value[1625] = 15'd3041;
    value[1626] = 15'd3045;
    value[1627] = 15'd3049;
    value[1628] = 15'd3053;
    value[1629] = 15'd3058;
    value[1630] = 15'd3062;
    value[1631] = 15'd3066;
    value[1632] = 15'd3070;
    value[1633] = 15'd3074;
    value[1634] = 15'd3078;
    value[1635] = 15'd3082;
    value[1636] = 15'd3086;
    value[1637] = 15'd3091;
    value[1638] = 15'd3095;
    value[1639] = 15'd3099;
    value[1640] = 15'd3103;
    value[1641] = 15'd3107;
    value[1642] = 15'd3111;
    value[1643] = 15'd3115;
    value[1644] = 15'd3119;
    value[1645] = 15'd3123;
    value[1646] = 15'd3128;
    value[1647] = 15'd3132;
    value[1648] = 15'd3136;
    value[1649] = 15'd3140;
    value[1650] = 15'd3144;
    value[1651] = 15'd3148;
    value[1652] = 15'd3152;
    value[1653] = 15'd3156;
    value[1654] = 15'd3160;
    value[1655] = 15'd3164;
    value[1656] = 15'd3168;
    value[1657] = 15'd3172;
    value[1658] = 15'd3176;
    value[1659] = 15'd3180;
    value[1660] = 15'd3184;
    value[1661] = 15'd3188;
    value[1662] = 15'd3192;
    value[1663] = 15'd3197;
    value[1664] = 15'd3201;
    value[1665] = 15'd3205;
    value[1666] = 15'd3209;
    value[1667] = 15'd3213;
    value[1668] = 15'd3217;
    value[1669] = 15'd3221;
    value[1670] = 15'd3225;
    value[1671] = 15'd3229;
    value[1672] = 15'd3233;
    value[1673] = 15'd3237;
    value[1674] = 15'd3241;
    value[1675] = 15'd3245;
    value[1676] = 15'd3249;
    value[1677] = 15'd3253;
    value[1678] = 15'd3257;
    value[1679] = 15'd3260;
    value[1680] = 15'd3264;
    value[1681] = 15'd3268;
    value[1682] = 15'd3272;
    value[1683] = 15'd3276;
    value[1684] = 15'd3280;
    value[1685] = 15'd3284;
    value[1686] = 15'd3288;
    value[1687] = 15'd3292;
    value[1688] = 15'd3296;
    value[1689] = 15'd3300;
    value[1690] = 15'd3304;
    value[1691] = 15'd3308;
    value[1692] = 15'd3312;
    value[1693] = 15'd3316;
    value[1694] = 15'd3320;
    value[1695] = 15'd3324;
    value[1696] = 15'd3327;
    value[1697] = 15'd3331;
    value[1698] = 15'd3335;
    value[1699] = 15'd3339;
    value[1700] = 15'd3343;
    value[1701] = 15'd3347;
    value[1702] = 15'd3351;
    value[1703] = 15'd3355;
    value[1704] = 15'd3359;
    value[1705] = 15'd3363;
    value[1706] = 15'd3366;
    value[1707] = 15'd3370;
    value[1708] = 15'd3374;
    value[1709] = 15'd3378;
    value[1710] = 15'd3382;
    value[1711] = 15'd3386;
    value[1712] = 15'd3390;
    value[1713] = 15'd3393;
    value[1714] = 15'd3397;
    value[1715] = 15'd3401;
    value[1716] = 15'd3405;
    value[1717] = 15'd3409;
    value[1718] = 15'd3413;
    value[1719] = 15'd3417;
    value[1720] = 15'd3420;
    value[1721] = 15'd3424;
    value[1722] = 15'd3428;
    value[1723] = 15'd3432;
    value[1724] = 15'd3436;
    value[1725] = 15'd3439;
    value[1726] = 15'd3443;
    value[1727] = 15'd3447;
    value[1728] = 15'd3451;
    value[1729] = 15'd3455;
    value[1730] = 15'd3458;
    value[1731] = 15'd3462;
    value[1732] = 15'd3466;
    value[1733] = 15'd3470;
    value[1734] = 15'd3474;
    value[1735] = 15'd3477;
    value[1736] = 15'd3481;
    value[1737] = 15'd3485;
    value[1738] = 15'd3489;
    value[1739] = 15'd3492;
    value[1740] = 15'd3496;
    value[1741] = 15'd3500;
    value[1742] = 15'd3504;
    value[1743] = 15'd3507;
    value[1744] = 15'd3511;
    value[1745] = 15'd3515;
    value[1746] = 15'd3519;
    value[1747] = 15'd3522;
    value[1748] = 15'd3526;
    value[1749] = 15'd3530;
    value[1750] = 15'd3534;
    value[1751] = 15'd3537;
    value[1752] = 15'd3541;
    value[1753] = 15'd3545;
    value[1754] = 15'd3548;
    value[1755] = 15'd3552;
    value[1756] = 15'd3556;
    value[1757] = 15'd3560;
    value[1758] = 15'd3563;
    value[1759] = 15'd3567;
    value[1760] = 15'd3571;
    value[1761] = 15'd3574;
    value[1762] = 15'd3578;
    value[1763] = 15'd3582;
    value[1764] = 15'd3585;
    value[1765] = 15'd3589;
    value[1766] = 15'd3593;
    value[1767] = 15'd3596;
    value[1768] = 15'd3600;
    value[1769] = 15'd3604;
    value[1770] = 15'd3607;
    value[1771] = 15'd3611;
    value[1772] = 15'd3615;
    value[1773] = 15'd3618;
    value[1774] = 15'd3622;
    value[1775] = 15'd3626;
    value[1776] = 15'd3629;
    value[1777] = 15'd3633;
    value[1778] = 15'd3637;
    value[1779] = 15'd3640;
    value[1780] = 15'd3644;
    value[1781] = 15'd3647;
    value[1782] = 15'd3651;
    value[1783] = 15'd3655;
    value[1784] = 15'd3658;
    value[1785] = 15'd3662;
    value[1786] = 15'd3665;
    value[1787] = 15'd3669;
    value[1788] = 15'd3673;
    value[1789] = 15'd3676;
    value[1790] = 15'd3680;
    value[1791] = 15'd3683;
    value[1792] = 15'd3687;
    value[1793] = 15'd3691;
    value[1794] = 15'd3694;
    value[1795] = 15'd3698;
    value[1796] = 15'd3701;
    value[1797] = 15'd3705;
    value[1798] = 15'd3708;
    value[1799] = 15'd3712;
    value[1800] = 15'd3716;
    value[1801] = 15'd3719;
    value[1802] = 15'd3723;
    value[1803] = 15'd3726;
    value[1804] = 15'd3730;
    value[1805] = 15'd3733;
    value[1806] = 15'd3737;
    value[1807] = 15'd3740;
    value[1808] = 15'd3744;
    value[1809] = 15'd3747;
    value[1810] = 15'd3751;
    value[1811] = 15'd3754;
    value[1812] = 15'd3758;
    value[1813] = 15'd3761;
    value[1814] = 15'd3765;
    value[1815] = 15'd3768;
    value[1816] = 15'd3772;
    value[1817] = 15'd3775;
    value[1818] = 15'd3779;
    value[1819] = 15'd3782;
    value[1820] = 15'd3786;
    value[1821] = 15'd3789;
    value[1822] = 15'd3793;
    value[1823] = 15'd3796;
    value[1824] = 15'd3800;
    value[1825] = 15'd3803;
    value[1826] = 15'd3807;
    value[1827] = 15'd3810;
    value[1828] = 15'd3814;
    value[1829] = 15'd3817;
    value[1830] = 15'd3821;
    value[1831] = 15'd3824;
    value[1832] = 15'd3828;
    value[1833] = 15'd3831;
    value[1834] = 15'd3834;
    value[1835] = 15'd3838;
    value[1836] = 15'd3841;
    value[1837] = 15'd3845;
    value[1838] = 15'd3848;
    value[1839] = 15'd3852;
    value[1840] = 15'd3855;
    value[1841] = 15'd3858;
    value[1842] = 15'd3862;
    value[1843] = 15'd3865;
    value[1844] = 15'd3869;
    value[1845] = 15'd3872;
    value[1846] = 15'd3876;
    value[1847] = 15'd3879;
    value[1848] = 15'd3882;
    value[1849] = 15'd3886;
    value[1850] = 15'd3889;
    value[1851] = 15'd3892;
    value[1852] = 15'd3896;
    value[1853] = 15'd3899;
    value[1854] = 15'd3903;
    value[1855] = 15'd3906;
    value[1856] = 15'd3909;
    value[1857] = 15'd3913;
    value[1858] = 15'd3916;
    value[1859] = 15'd3919;
    value[1860] = 15'd3923;
    value[1861] = 15'd3926;
    value[1862] = 15'd3930;
    value[1863] = 15'd3933;
    value[1864] = 15'd3936;
    value[1865] = 15'd3940;
    value[1866] = 15'd3943;
    value[1867] = 15'd3946;
    value[1868] = 15'd3950;
    value[1869] = 15'd3953;
    value[1870] = 15'd3956;
    value[1871] = 15'd3960;
    value[1872] = 15'd3963;
    value[1873] = 15'd3966;
    value[1874] = 15'd3970;
    value[1875] = 15'd3973;
    value[1876] = 15'd3976;
    value[1877] = 15'd3979;
    value[1878] = 15'd3983;
    value[1879] = 15'd3986;
    value[1880] = 15'd3989;
    value[1881] = 15'd3993;
    value[1882] = 15'd3996;
    value[1883] = 15'd3999;
    value[1884] = 15'd4003;
    value[1885] = 15'd4006;
    value[1886] = 15'd4009;
    value[1887] = 15'd4012;
    value[1888] = 15'd4016;
    value[1889] = 15'd4019;
    value[1890] = 15'd4022;
    value[1891] = 15'd4025;
    value[1892] = 15'd4029;
    value[1893] = 15'd4032;
    value[1894] = 15'd4035;
    value[1895] = 15'd4038;
    value[1896] = 15'd4042;
    value[1897] = 15'd4045;
    value[1898] = 15'd4048;
    value[1899] = 15'd4051;
    value[1900] = 15'd4055;
    value[1901] = 15'd4058;
    value[1902] = 15'd4061;
    value[1903] = 15'd4064;
    value[1904] = 15'd4067;
    value[1905] = 15'd4071;
    value[1906] = 15'd4074;
    value[1907] = 15'd4077;
    value[1908] = 15'd4080;
    value[1909] = 15'd4084;
    value[1910] = 15'd4087;
    value[1911] = 15'd4090;
    value[1912] = 15'd4093;
    value[1913] = 15'd4096;
    value[1914] = 15'd4100;
    value[1915] = 15'd4103;
    value[1916] = 15'd4106;
    value[1917] = 15'd4109;
    value[1918] = 15'd4112;
    value[1919] = 15'd4115;
    value[1920] = 15'd4119;
    value[1921] = 15'd4122;
    value[1922] = 15'd4125;
    value[1923] = 15'd4128;
    value[1924] = 15'd4131;
    value[1925] = 15'd4134;
    value[1926] = 15'd4138;
    value[1927] = 15'd4141;
    value[1928] = 15'd4144;
    value[1929] = 15'd4147;
    value[1930] = 15'd4150;
    value[1931] = 15'd4153;
    value[1932] = 15'd4156;
    value[1933] = 15'd4160;
    value[1934] = 15'd4163;
    value[1935] = 15'd4166;
    value[1936] = 15'd4169;
    value[1937] = 15'd4172;
    value[1938] = 15'd4175;
    value[1939] = 15'd4178;
    value[1940] = 15'd4181;
    value[1941] = 15'd4184;
    value[1942] = 15'd4188;
    value[1943] = 15'd4191;
    value[1944] = 15'd4194;
    value[1945] = 15'd4197;
    value[1946] = 15'd4200;
    value[1947] = 15'd4203;
    value[1948] = 15'd4206;
    value[1949] = 15'd4209;
    value[1950] = 15'd4212;
    value[1951] = 15'd4215;
    value[1952] = 15'd4218;
    value[1953] = 15'd4222;
    value[1954] = 15'd4225;
    value[1955] = 15'd4228;
    value[1956] = 15'd4231;
    value[1957] = 15'd4234;
    value[1958] = 15'd4237;
    value[1959] = 15'd4240;
    value[1960] = 15'd4243;
    value[1961] = 15'd4246;
    value[1962] = 15'd4249;
    value[1963] = 15'd4252;
    value[1964] = 15'd4255;
    value[1965] = 15'd4258;
    value[1966] = 15'd4261;
    value[1967] = 15'd4264;
    value[1968] = 15'd4267;
    value[1969] = 15'd4270;
    value[1970] = 15'd4273;
    value[1971] = 15'd4276;
    value[1972] = 15'd4279;
    value[1973] = 15'd4282;
    value[1974] = 15'd4285;
    value[1975] = 15'd4288;
    value[1976] = 15'd4291;
    value[1977] = 15'd4294;
    value[1978] = 15'd4297;
    value[1979] = 15'd4300;
    value[1980] = 15'd4303;
    value[1981] = 15'd4306;
    value[1982] = 15'd4309;
    value[1983] = 15'd4312;
    value[1984] = 15'd4315;
    value[1985] = 15'd4318;
    value[1986] = 15'd4321;
    value[1987] = 15'd4324;
    value[1988] = 15'd4327;
    value[1989] = 15'd4330;
    value[1990] = 15'd4333;
    value[1991] = 15'd4336;
    value[1992] = 15'd4339;
    value[1993] = 15'd4342;
    value[1994] = 15'd4345;
    value[1995] = 15'd4348;
    value[1996] = 15'd4351;
    value[1997] = 15'd4354;
    value[1998] = 15'd4357;
    value[1999] = 15'd4360;
    value[2000] = 15'd4363;
    value[2001] = 15'd4365;
    value[2002] = 15'd4368;
    value[2003] = 15'd4371;
    value[2004] = 15'd4374;
    value[2005] = 15'd4377;
    value[2006] = 15'd4380;
    value[2007] = 15'd4383;
    value[2008] = 15'd4386;
    value[2009] = 15'd4389;
    value[2010] = 15'd4392;
    value[2011] = 15'd4395;
    value[2012] = 15'd4397;
    value[2013] = 15'd4400;
    value[2014] = 15'd4403;
    value[2015] = 15'd4406;
    value[2016] = 15'd4409;
    value[2017] = 15'd4412;
    value[2018] = 15'd4415;
    value[2019] = 15'd4418;
    value[2020] = 15'd4421;
    value[2021] = 15'd4423;
    value[2022] = 15'd4426;
    value[2023] = 15'd4429;
    value[2024] = 15'd4432;
    value[2025] = 15'd4435;
    value[2026] = 15'd4438;
    value[2027] = 15'd4441;
    value[2028] = 15'd4443;
    value[2029] = 15'd4446;
    value[2030] = 15'd4449;
    value[2031] = 15'd4452;
    value[2032] = 15'd4455;
    value[2033] = 15'd4458;
    value[2034] = 15'd4461;
    value[2035] = 15'd4463;
    value[2036] = 15'd4466;
    value[2037] = 15'd4469;
    value[2038] = 15'd4472;
    value[2039] = 15'd4475;
    value[2040] = 15'd4478;
    value[2041] = 15'd4480;
    value[2042] = 15'd4483;
    value[2043] = 15'd4486;
    value[2044] = 15'd4489;
    value[2045] = 15'd4492;
    value[2046] = 15'd4494;
    value[2047] = 15'd4497;

  end

endmodule
