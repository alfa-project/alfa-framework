/*
 * Copyright 2025 ALFA Project. All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`timescale 1ns / 1ps

module alib_cos (
    input i_clk,
    input i_rst,
    input [15:0] i_angle,
    output wire [16:0] o_value,
    output wire [0:0] o_sig
);

  wire [15:0] true_angle;
  wire [16:0] value      [9000:0];

  assign true_angle = i_angle > 35999 ? i_angle - 35999 : i_angle;

  assign true_angle = i_angle > 35999 ? i_angle - 35999 : i_angle;

  assign o_value = (true_angle>0 && true_angle<9000) ? value[true_angle] : 
                   (true_angle>9000 && true_angle<18000) ? value[18000-true_angle] : 
                   (true_angle>18000 && true_angle<27000) ? value[true_angle-18000] : 
                   value[36000-true_angle];

  assign o_sig = ((i_angle < 9001) || (i_angle > 27000)) ? 0 : 1;

  initial begin

    value[0] = 17'd100000;
    value[1] = 17'd100000;
    value[2] = 17'd99999;
    value[3] = 17'd99999;
    value[4] = 17'd99999;
    value[5] = 17'd99999;
    value[6] = 17'd99999;
    value[7] = 17'd99999;
    value[8] = 17'd99999;
    value[9] = 17'd99999;
    value[10] = 17'd99999;
    value[11] = 17'd99999;
    value[12] = 17'd99999;
    value[13] = 17'd99999;
    value[14] = 17'd99999;
    value[15] = 17'd99999;
    value[16] = 17'd99999;
    value[17] = 17'd99999;
    value[18] = 17'd99999;
    value[19] = 17'd99999;
    value[20] = 17'd99999;
    value[21] = 17'd99999;
    value[22] = 17'd99999;
    value[23] = 17'd99999;
    value[24] = 17'd99999;
    value[25] = 17'd99999;
    value[26] = 17'd99998;
    value[27] = 17'd99998;
    value[28] = 17'd99998;
    value[29] = 17'd99998;
    value[30] = 17'd99998;
    value[31] = 17'd99998;
    value[32] = 17'd99998;
    value[33] = 17'd99998;
    value[34] = 17'd99998;
    value[35] = 17'd99998;
    value[36] = 17'd99998;
    value[37] = 17'd99997;
    value[38] = 17'd99997;
    value[39] = 17'd99997;
    value[40] = 17'd99997;
    value[41] = 17'd99997;
    value[42] = 17'd99997;
    value[43] = 17'd99997;
    value[44] = 17'd99997;
    value[45] = 17'd99996;
    value[46] = 17'd99996;
    value[47] = 17'd99996;
    value[48] = 17'd99996;
    value[49] = 17'd99996;
    value[50] = 17'd99996;
    value[51] = 17'd99996;
    value[52] = 17'd99995;
    value[53] = 17'd99995;
    value[54] = 17'd99995;
    value[55] = 17'd99995;
    value[56] = 17'd99995;
    value[57] = 17'd99995;
    value[58] = 17'd99994;
    value[59] = 17'd99994;
    value[60] = 17'd99994;
    value[61] = 17'd99994;
    value[62] = 17'd99994;
    value[63] = 17'd99993;
    value[64] = 17'd99993;
    value[65] = 17'd99993;
    value[66] = 17'd99993;
    value[67] = 17'd99993;
    value[68] = 17'd99992;
    value[69] = 17'd99992;
    value[70] = 17'd99992;
    value[71] = 17'd99992;
    value[72] = 17'd99992;
    value[73] = 17'd99991;
    value[74] = 17'd99991;
    value[75] = 17'd99991;
    value[76] = 17'd99991;
    value[77] = 17'd99990;
    value[78] = 17'd99990;
    value[79] = 17'd99990;
    value[80] = 17'd99990;
    value[81] = 17'd99990;
    value[82] = 17'd99989;
    value[83] = 17'd99989;
    value[84] = 17'd99989;
    value[85] = 17'd99988;
    value[86] = 17'd99988;
    value[87] = 17'd99988;
    value[88] = 17'd99988;
    value[89] = 17'd99987;
    value[90] = 17'd99987;
    value[91] = 17'd99987;
    value[92] = 17'd99987;
    value[93] = 17'd99986;
    value[94] = 17'd99986;
    value[95] = 17'd99986;
    value[96] = 17'd99985;
    value[97] = 17'd99985;
    value[98] = 17'd99985;
    value[99] = 17'd99985;
    value[100] = 17'd99984;
    value[101] = 17'd99984;
    value[102] = 17'd99984;
    value[103] = 17'd99983;
    value[104] = 17'd99983;
    value[105] = 17'd99983;
    value[106] = 17'd99982;
    value[107] = 17'd99982;
    value[108] = 17'd99982;
    value[109] = 17'd99981;
    value[110] = 17'd99981;
    value[111] = 17'd99981;
    value[112] = 17'd99980;
    value[113] = 17'd99980;
    value[114] = 17'd99980;
    value[115] = 17'd99979;
    value[116] = 17'd99979;
    value[117] = 17'd99979;
    value[118] = 17'd99978;
    value[119] = 17'd99978;
    value[120] = 17'd99978;
    value[121] = 17'd99977;
    value[122] = 17'd99977;
    value[123] = 17'd99976;
    value[124] = 17'd99976;
    value[125] = 17'd99976;
    value[126] = 17'd99975;
    value[127] = 17'd99975;
    value[128] = 17'd99975;
    value[129] = 17'd99974;
    value[130] = 17'd99974;
    value[131] = 17'd99973;
    value[132] = 17'd99973;
    value[133] = 17'd99973;
    value[134] = 17'd99972;
    value[135] = 17'd99972;
    value[136] = 17'd99971;
    value[137] = 17'd99971;
    value[138] = 17'd99970;
    value[139] = 17'd99970;
    value[140] = 17'd99970;
    value[141] = 17'd99969;
    value[142] = 17'd99969;
    value[143] = 17'd99968;
    value[144] = 17'd99968;
    value[145] = 17'd99967;
    value[146] = 17'd99967;
    value[147] = 17'd99967;
    value[148] = 17'd99966;
    value[149] = 17'd99966;
    value[150] = 17'd99965;
    value[151] = 17'd99965;
    value[152] = 17'd99964;
    value[153] = 17'd99964;
    value[154] = 17'd99963;
    value[155] = 17'd99963;
    value[156] = 17'd99962;
    value[157] = 17'd99962;
    value[158] = 17'd99961;
    value[159] = 17'd99961;
    value[160] = 17'd99961;
    value[161] = 17'd99960;
    value[162] = 17'd99960;
    value[163] = 17'd99959;
    value[164] = 17'd99959;
    value[165] = 17'd99958;
    value[166] = 17'd99958;
    value[167] = 17'd99957;
    value[168] = 17'd99957;
    value[169] = 17'd99956;
    value[170] = 17'd99955;
    value[171] = 17'd99955;
    value[172] = 17'd99954;
    value[173] = 17'd99954;
    value[174] = 17'd99953;
    value[175] = 17'd99953;
    value[176] = 17'd99952;
    value[177] = 17'd99952;
    value[178] = 17'd99951;
    value[179] = 17'd99951;
    value[180] = 17'd99950;
    value[181] = 17'd99950;
    value[182] = 17'd99949;
    value[183] = 17'd99949;
    value[184] = 17'd99948;
    value[185] = 17'd99947;
    value[186] = 17'd99947;
    value[187] = 17'd99946;
    value[188] = 17'd99946;
    value[189] = 17'd99945;
    value[190] = 17'd99945;
    value[191] = 17'd99944;
    value[192] = 17'd99943;
    value[193] = 17'd99943;
    value[194] = 17'd99942;
    value[195] = 17'd99942;
    value[196] = 17'd99941;
    value[197] = 17'd99940;
    value[198] = 17'd99940;
    value[199] = 17'd99939;
    value[200] = 17'd99939;
    value[201] = 17'd99938;
    value[202] = 17'd99937;
    value[203] = 17'd99937;
    value[204] = 17'd99936;
    value[205] = 17'd99936;
    value[206] = 17'd99935;
    value[207] = 17'd99934;
    value[208] = 17'd99934;
    value[209] = 17'd99933;
    value[210] = 17'd99932;
    value[211] = 17'd99932;
    value[212] = 17'd99931;
    value[213] = 17'd99930;
    value[214] = 17'd99930;
    value[215] = 17'd99929;
    value[216] = 17'd99928;
    value[217] = 17'd99928;
    value[218] = 17'd99927;
    value[219] = 17'd99926;
    value[220] = 17'd99926;
    value[221] = 17'd99925;
    value[222] = 17'd99924;
    value[223] = 17'd99924;
    value[224] = 17'd99923;
    value[225] = 17'd99922;
    value[226] = 17'd99922;
    value[227] = 17'd99921;
    value[228] = 17'd99920;
    value[229] = 17'd99920;
    value[230] = 17'd99919;
    value[231] = 17'd99918;
    value[232] = 17'd99918;
    value[233] = 17'd99917;
    value[234] = 17'd99916;
    value[235] = 17'd99915;
    value[236] = 17'd99915;
    value[237] = 17'd99914;
    value[238] = 17'd99913;
    value[239] = 17'd99913;
    value[240] = 17'd99912;
    value[241] = 17'd99911;
    value[242] = 17'd99910;
    value[243] = 17'd99910;
    value[244] = 17'd99909;
    value[245] = 17'd99908;
    value[246] = 17'd99907;
    value[247] = 17'd99907;
    value[248] = 17'd99906;
    value[249] = 17'd99905;
    value[250] = 17'd99904;
    value[251] = 17'd99904;
    value[252] = 17'd99903;
    value[253] = 17'd99902;
    value[254] = 17'd99901;
    value[255] = 17'd99900;
    value[256] = 17'd99900;
    value[257] = 17'd99899;
    value[258] = 17'd99898;
    value[259] = 17'd99897;
    value[260] = 17'd99897;
    value[261] = 17'd99896;
    value[262] = 17'd99895;
    value[263] = 17'd99894;
    value[264] = 17'd99893;
    value[265] = 17'd99893;
    value[266] = 17'd99892;
    value[267] = 17'd99891;
    value[268] = 17'd99890;
    value[269] = 17'd99889;
    value[270] = 17'd99888;
    value[271] = 17'd99888;
    value[272] = 17'd99887;
    value[273] = 17'd99886;
    value[274] = 17'd99885;
    value[275] = 17'd99884;
    value[276] = 17'd99884;
    value[277] = 17'd99883;
    value[278] = 17'd99882;
    value[279] = 17'd99881;
    value[280] = 17'd99880;
    value[281] = 17'd99879;
    value[282] = 17'd99878;
    value[283] = 17'd99878;
    value[284] = 17'd99877;
    value[285] = 17'd99876;
    value[286] = 17'd99875;
    value[287] = 17'd99874;
    value[288] = 17'd99873;
    value[289] = 17'd99872;
    value[290] = 17'd99871;
    value[291] = 17'd99871;
    value[292] = 17'd99870;
    value[293] = 17'd99869;
    value[294] = 17'd99868;
    value[295] = 17'd99867;
    value[296] = 17'd99866;
    value[297] = 17'd99865;
    value[298] = 17'd99864;
    value[299] = 17'd99863;
    value[300] = 17'd99862;
    value[301] = 17'd99862;
    value[302] = 17'd99861;
    value[303] = 17'd99860;
    value[304] = 17'd99859;
    value[305] = 17'd99858;
    value[306] = 17'd99857;
    value[307] = 17'd99856;
    value[308] = 17'd99855;
    value[309] = 17'd99854;
    value[310] = 17'd99853;
    value[311] = 17'd99852;
    value[312] = 17'd99851;
    value[313] = 17'd99850;
    value[314] = 17'd99849;
    value[315] = 17'd99848;
    value[316] = 17'd99847;
    value[317] = 17'd99846;
    value[318] = 17'd99846;
    value[319] = 17'd99845;
    value[320] = 17'd99844;
    value[321] = 17'd99843;
    value[322] = 17'd99842;
    value[323] = 17'd99841;
    value[324] = 17'd99840;
    value[325] = 17'd99839;
    value[326] = 17'd99838;
    value[327] = 17'd99837;
    value[328] = 17'd99836;
    value[329] = 17'd99835;
    value[330] = 17'd99834;
    value[331] = 17'd99833;
    value[332] = 17'd99832;
    value[333] = 17'd99831;
    value[334] = 17'd99830;
    value[335] = 17'd99829;
    value[336] = 17'd99828;
    value[337] = 17'd99827;
    value[338] = 17'd99826;
    value[339] = 17'd99825;
    value[340] = 17'd99823;
    value[341] = 17'd99822;
    value[342] = 17'd99821;
    value[343] = 17'd99820;
    value[344] = 17'd99819;
    value[345] = 17'd99818;
    value[346] = 17'd99817;
    value[347] = 17'd99816;
    value[348] = 17'd99815;
    value[349] = 17'd99814;
    value[350] = 17'd99813;
    value[351] = 17'd99812;
    value[352] = 17'd99811;
    value[353] = 17'd99810;
    value[354] = 17'd99809;
    value[355] = 17'd99808;
    value[356] = 17'd99807;
    value[357] = 17'd99805;
    value[358] = 17'd99804;
    value[359] = 17'd99803;
    value[360] = 17'd99802;
    value[361] = 17'd99801;
    value[362] = 17'd99800;
    value[363] = 17'd99799;
    value[364] = 17'd99798;
    value[365] = 17'd99797;
    value[366] = 17'd99796;
    value[367] = 17'd99794;
    value[368] = 17'd99793;
    value[369] = 17'd99792;
    value[370] = 17'd99791;
    value[371] = 17'd99790;
    value[372] = 17'd99789;
    value[373] = 17'd99788;
    value[374] = 17'd99787;
    value[375] = 17'd99785;
    value[376] = 17'd99784;
    value[377] = 17'd99783;
    value[378] = 17'd99782;
    value[379] = 17'd99781;
    value[380] = 17'd99780;
    value[381] = 17'd99778;
    value[382] = 17'd99777;
    value[383] = 17'd99776;
    value[384] = 17'd99775;
    value[385] = 17'd99774;
    value[386] = 17'd99773;
    value[387] = 17'd99771;
    value[388] = 17'd99770;
    value[389] = 17'd99769;
    value[390] = 17'd99768;
    value[391] = 17'd99767;
    value[392] = 17'd99766;
    value[393] = 17'd99764;
    value[394] = 17'd99763;
    value[395] = 17'd99762;
    value[396] = 17'd99761;
    value[397] = 17'd99760;
    value[398] = 17'd99758;
    value[399] = 17'd99757;
    value[400] = 17'd99756;
    value[401] = 17'd99755;
    value[402] = 17'd99753;
    value[403] = 17'd99752;
    value[404] = 17'd99751;
    value[405] = 17'd99750;
    value[406] = 17'd99749;
    value[407] = 17'd99747;
    value[408] = 17'd99746;
    value[409] = 17'd99745;
    value[410] = 17'd99744;
    value[411] = 17'd99742;
    value[412] = 17'd99741;
    value[413] = 17'd99740;
    value[414] = 17'd99739;
    value[415] = 17'd99737;
    value[416] = 17'd99736;
    value[417] = 17'd99735;
    value[418] = 17'd99734;
    value[419] = 17'd99732;
    value[420] = 17'd99731;
    value[421] = 17'd99730;
    value[422] = 17'd99728;
    value[423] = 17'd99727;
    value[424] = 17'd99726;
    value[425] = 17'd99725;
    value[426] = 17'd99723;
    value[427] = 17'd99722;
    value[428] = 17'd99721;
    value[429] = 17'd99719;
    value[430] = 17'd99718;
    value[431] = 17'd99717;
    value[432] = 17'd99715;
    value[433] = 17'd99714;
    value[434] = 17'd99713;
    value[435] = 17'd99711;
    value[436] = 17'd99710;
    value[437] = 17'd99709;
    value[438] = 17'd99707;
    value[439] = 17'd99706;
    value[440] = 17'd99705;
    value[441] = 17'd99703;
    value[442] = 17'd99702;
    value[443] = 17'd99701;
    value[444] = 17'd99699;
    value[445] = 17'd99698;
    value[446] = 17'd99697;
    value[447] = 17'd99695;
    value[448] = 17'd99694;
    value[449] = 17'd99693;
    value[450] = 17'd99691;
    value[451] = 17'd99690;
    value[452] = 17'd99688;
    value[453] = 17'd99687;
    value[454] = 17'd99686;
    value[455] = 17'd99684;
    value[456] = 17'd99683;
    value[457] = 17'd99682;
    value[458] = 17'd99680;
    value[459] = 17'd99679;
    value[460] = 17'd99677;
    value[461] = 17'd99676;
    value[462] = 17'd99675;
    value[463] = 17'd99673;
    value[464] = 17'd99672;
    value[465] = 17'd99670;
    value[466] = 17'd99669;
    value[467] = 17'd99668;
    value[468] = 17'd99666;
    value[469] = 17'd99665;
    value[470] = 17'd99663;
    value[471] = 17'd99662;
    value[472] = 17'd99660;
    value[473] = 17'd99659;
    value[474] = 17'd99657;
    value[475] = 17'd99656;
    value[476] = 17'd99655;
    value[477] = 17'd99653;
    value[478] = 17'd99652;
    value[479] = 17'd99650;
    value[480] = 17'd99649;
    value[481] = 17'd99647;
    value[482] = 17'd99646;
    value[483] = 17'd99644;
    value[484] = 17'd99643;
    value[485] = 17'd99641;
    value[486] = 17'd99640;
    value[487] = 17'd99638;
    value[488] = 17'd99637;
    value[489] = 17'd99636;
    value[490] = 17'd99634;
    value[491] = 17'd99633;
    value[492] = 17'd99631;
    value[493] = 17'd99630;
    value[494] = 17'd99628;
    value[495] = 17'd99627;
    value[496] = 17'd99625;
    value[497] = 17'd99624;
    value[498] = 17'd99622;
    value[499] = 17'd99620;
    value[500] = 17'd99619;
    value[501] = 17'd99617;
    value[502] = 17'd99616;
    value[503] = 17'd99614;
    value[504] = 17'd99613;
    value[505] = 17'd99611;
    value[506] = 17'd99610;
    value[507] = 17'd99608;
    value[508] = 17'd99607;
    value[509] = 17'd99605;
    value[510] = 17'd99604;
    value[511] = 17'd99602;
    value[512] = 17'd99601;
    value[513] = 17'd99599;
    value[514] = 17'd99597;
    value[515] = 17'd99596;
    value[516] = 17'd99594;
    value[517] = 17'd99593;
    value[518] = 17'd99591;
    value[519] = 17'd99590;
    value[520] = 17'd99588;
    value[521] = 17'd99586;
    value[522] = 17'd99585;
    value[523] = 17'd99583;
    value[524] = 17'd99582;
    value[525] = 17'd99580;
    value[526] = 17'd99578;
    value[527] = 17'd99577;
    value[528] = 17'd99575;
    value[529] = 17'd99574;
    value[530] = 17'd99572;
    value[531] = 17'd99570;
    value[532] = 17'd99569;
    value[533] = 17'd99567;
    value[534] = 17'd99566;
    value[535] = 17'd99564;
    value[536] = 17'd99562;
    value[537] = 17'd99561;
    value[538] = 17'd99559;
    value[539] = 17'd99557;
    value[540] = 17'd99556;
    value[541] = 17'd99554;
    value[542] = 17'd99552;
    value[543] = 17'd99551;
    value[544] = 17'd99549;
    value[545] = 17'd99547;
    value[546] = 17'd99546;
    value[547] = 17'd99544;
    value[548] = 17'd99542;
    value[549] = 17'd99541;
    value[550] = 17'd99539;
    value[551] = 17'd99537;
    value[552] = 17'd99536;
    value[553] = 17'd99534;
    value[554] = 17'd99532;
    value[555] = 17'd99531;
    value[556] = 17'd99529;
    value[557] = 17'd99527;
    value[558] = 17'd99526;
    value[559] = 17'd99524;
    value[560] = 17'd99522;
    value[561] = 17'd99521;
    value[562] = 17'd99519;
    value[563] = 17'd99517;
    value[564] = 17'd99515;
    value[565] = 17'd99514;
    value[566] = 17'd99512;
    value[567] = 17'd99510;
    value[568] = 17'd99509;
    value[569] = 17'd99507;
    value[570] = 17'd99505;
    value[571] = 17'd99503;
    value[572] = 17'd99502;
    value[573] = 17'd99500;
    value[574] = 17'd99498;
    value[575] = 17'd99496;
    value[576] = 17'd99495;
    value[577] = 17'd99493;
    value[578] = 17'd99491;
    value[579] = 17'd99489;
    value[580] = 17'd99488;
    value[581] = 17'd99486;
    value[582] = 17'd99484;
    value[583] = 17'd99482;
    value[584] = 17'd99480;
    value[585] = 17'd99479;
    value[586] = 17'd99477;
    value[587] = 17'd99475;
    value[588] = 17'd99473;
    value[589] = 17'd99472;
    value[590] = 17'd99470;
    value[591] = 17'd99468;
    value[592] = 17'd99466;
    value[593] = 17'd99464;
    value[594] = 17'd99463;
    value[595] = 17'd99461;
    value[596] = 17'd99459;
    value[597] = 17'd99457;
    value[598] = 17'd99455;
    value[599] = 17'd99454;
    value[600] = 17'd99452;
    value[601] = 17'd99450;
    value[602] = 17'd99448;
    value[603] = 17'd99446;
    value[604] = 17'd99444;
    value[605] = 17'd99443;
    value[606] = 17'd99441;
    value[607] = 17'd99439;
    value[608] = 17'd99437;
    value[609] = 17'd99435;
    value[610] = 17'd99433;
    value[611] = 17'd99431;
    value[612] = 17'd99430;
    value[613] = 17'd99428;
    value[614] = 17'd99426;
    value[615] = 17'd99424;
    value[616] = 17'd99422;
    value[617] = 17'd99420;
    value[618] = 17'd99418;
    value[619] = 17'd99416;
    value[620] = 17'd99415;
    value[621] = 17'd99413;
    value[622] = 17'd99411;
    value[623] = 17'd99409;
    value[624] = 17'd99407;
    value[625] = 17'd99405;
    value[626] = 17'd99403;
    value[627] = 17'd99401;
    value[628] = 17'd99399;
    value[629] = 17'd99398;
    value[630] = 17'd99396;
    value[631] = 17'd99394;
    value[632] = 17'd99392;
    value[633] = 17'd99390;
    value[634] = 17'd99388;
    value[635] = 17'd99386;
    value[636] = 17'd99384;
    value[637] = 17'd99382;
    value[638] = 17'd99380;
    value[639] = 17'd99378;
    value[640] = 17'd99376;
    value[641] = 17'd99374;
    value[642] = 17'd99372;
    value[643] = 17'd99370;
    value[644] = 17'd99368;
    value[645] = 17'd99367;
    value[646] = 17'd99365;
    value[647] = 17'd99363;
    value[648] = 17'd99361;
    value[649] = 17'd99359;
    value[650] = 17'd99357;
    value[651] = 17'd99355;
    value[652] = 17'd99353;
    value[653] = 17'd99351;
    value[654] = 17'd99349;
    value[655] = 17'd99347;
    value[656] = 17'd99345;
    value[657] = 17'd99343;
    value[658] = 17'd99341;
    value[659] = 17'd99339;
    value[660] = 17'd99337;
    value[661] = 17'd99335;
    value[662] = 17'd99333;
    value[663] = 17'd99331;
    value[664] = 17'd99329;
    value[665] = 17'd99327;
    value[666] = 17'd99325;
    value[667] = 17'd99323;
    value[668] = 17'd99321;
    value[669] = 17'd99319;
    value[670] = 17'd99317;
    value[671] = 17'd99315;
    value[672] = 17'd99312;
    value[673] = 17'd99310;
    value[674] = 17'd99308;
    value[675] = 17'd99306;
    value[676] = 17'd99304;
    value[677] = 17'd99302;
    value[678] = 17'd99300;
    value[679] = 17'd99298;
    value[680] = 17'd99296;
    value[681] = 17'd99294;
    value[682] = 17'd99292;
    value[683] = 17'd99290;
    value[684] = 17'd99288;
    value[685] = 17'd99286;
    value[686] = 17'd99284;
    value[687] = 17'd99282;
    value[688] = 17'd99279;
    value[689] = 17'd99277;
    value[690] = 17'd99275;
    value[691] = 17'd99273;
    value[692] = 17'd99271;
    value[693] = 17'd99269;
    value[694] = 17'd99267;
    value[695] = 17'd99265;
    value[696] = 17'd99263;
    value[697] = 17'd99260;
    value[698] = 17'd99258;
    value[699] = 17'd99256;
    value[700] = 17'd99254;
    value[701] = 17'd99252;
    value[702] = 17'd99250;
    value[703] = 17'd99248;
    value[704] = 17'd99246;
    value[705] = 17'd99243;
    value[706] = 17'd99241;
    value[707] = 17'd99239;
    value[708] = 17'd99237;
    value[709] = 17'd99235;
    value[710] = 17'd99233;
    value[711] = 17'd99231;
    value[712] = 17'd99228;
    value[713] = 17'd99226;
    value[714] = 17'd99224;
    value[715] = 17'd99222;
    value[716] = 17'd99220;
    value[717] = 17'd99218;
    value[718] = 17'd99215;
    value[719] = 17'd99213;
    value[720] = 17'd99211;
    value[721] = 17'd99209;
    value[722] = 17'd99207;
    value[723] = 17'd99204;
    value[724] = 17'd99202;
    value[725] = 17'd99200;
    value[726] = 17'd99198;
    value[727] = 17'd99196;
    value[728] = 17'd99193;
    value[729] = 17'd99191;
    value[730] = 17'd99189;
    value[731] = 17'd99187;
    value[732] = 17'd99185;
    value[733] = 17'd99182;
    value[734] = 17'd99180;
    value[735] = 17'd99178;
    value[736] = 17'd99176;
    value[737] = 17'd99173;
    value[738] = 17'd99171;
    value[739] = 17'd99169;
    value[740] = 17'd99167;
    value[741] = 17'd99164;
    value[742] = 17'd99162;
    value[743] = 17'd99160;
    value[744] = 17'd99158;
    value[745] = 17'd99155;
    value[746] = 17'd99153;
    value[747] = 17'd99151;
    value[748] = 17'd99149;
    value[749] = 17'd99146;
    value[750] = 17'd99144;
    value[751] = 17'd99142;
    value[752] = 17'd99139;
    value[753] = 17'd99137;
    value[754] = 17'd99135;
    value[755] = 17'd99133;
    value[756] = 17'd99130;
    value[757] = 17'd99128;
    value[758] = 17'd99126;
    value[759] = 17'd99123;
    value[760] = 17'd99121;
    value[761] = 17'd99119;
    value[762] = 17'd99116;
    value[763] = 17'd99114;
    value[764] = 17'd99112;
    value[765] = 17'd99109;
    value[766] = 17'd99107;
    value[767] = 17'd99105;
    value[768] = 17'd99102;
    value[769] = 17'd99100;
    value[770] = 17'd99098;
    value[771] = 17'd99095;
    value[772] = 17'd99093;
    value[773] = 17'd99091;
    value[774] = 17'd99088;
    value[775] = 17'd99086;
    value[776] = 17'd99084;
    value[777] = 17'd99081;
    value[778] = 17'd99079;
    value[779] = 17'd99077;
    value[780] = 17'd99074;
    value[781] = 17'd99072;
    value[782] = 17'd99070;
    value[783] = 17'd99067;
    value[784] = 17'd99065;
    value[785] = 17'd99062;
    value[786] = 17'd99060;
    value[787] = 17'd99058;
    value[788] = 17'd99055;
    value[789] = 17'd99053;
    value[790] = 17'd99050;
    value[791] = 17'd99048;
    value[792] = 17'd99046;
    value[793] = 17'd99043;
    value[794] = 17'd99041;
    value[795] = 17'd99038;
    value[796] = 17'd99036;
    value[797] = 17'd99034;
    value[798] = 17'd99031;
    value[799] = 17'd99029;
    value[800] = 17'd99026;
    value[801] = 17'd99024;
    value[802] = 17'd99021;
    value[803] = 17'd99019;
    value[804] = 17'd99017;
    value[805] = 17'd99014;
    value[806] = 17'd99012;
    value[807] = 17'd99009;
    value[808] = 17'd99007;
    value[809] = 17'd99004;
    value[810] = 17'd99002;
    value[811] = 17'd98999;
    value[812] = 17'd98997;
    value[813] = 17'd98994;
    value[814] = 17'd98992;
    value[815] = 17'd98990;
    value[816] = 17'd98987;
    value[817] = 17'd98985;
    value[818] = 17'd98982;
    value[819] = 17'd98980;
    value[820] = 17'd98977;
    value[821] = 17'd98975;
    value[822] = 17'd98972;
    value[823] = 17'd98970;
    value[824] = 17'd98967;
    value[825] = 17'd98965;
    value[826] = 17'd98962;
    value[827] = 17'd98960;
    value[828] = 17'd98957;
    value[829] = 17'd98955;
    value[830] = 17'd98952;
    value[831] = 17'd98950;
    value[832] = 17'd98947;
    value[833] = 17'd98945;
    value[834] = 17'd98942;
    value[835] = 17'd98939;
    value[836] = 17'd98937;
    value[837] = 17'd98934;
    value[838] = 17'd98932;
    value[839] = 17'd98929;
    value[840] = 17'd98927;
    value[841] = 17'd98924;
    value[842] = 17'd98922;
    value[843] = 17'd98919;
    value[844] = 17'd98917;
    value[845] = 17'd98914;
    value[846] = 17'd98911;
    value[847] = 17'd98909;
    value[848] = 17'd98906;
    value[849] = 17'd98904;
    value[850] = 17'd98901;
    value[851] = 17'd98899;
    value[852] = 17'd98896;
    value[853] = 17'd98893;
    value[854] = 17'd98891;
    value[855] = 17'd98888;
    value[856] = 17'd98886;
    value[857] = 17'd98883;
    value[858] = 17'd98880;
    value[859] = 17'd98878;
    value[860] = 17'd98875;
    value[861] = 17'd98873;
    value[862] = 17'd98870;
    value[863] = 17'd98867;
    value[864] = 17'd98865;
    value[865] = 17'd98862;
    value[866] = 17'd98859;
    value[867] = 17'd98857;
    value[868] = 17'd98854;
    value[869] = 17'd98852;
    value[870] = 17'd98849;
    value[871] = 17'd98846;
    value[872] = 17'd98844;
    value[873] = 17'd98841;
    value[874] = 17'd98838;
    value[875] = 17'd98836;
    value[876] = 17'd98833;
    value[877] = 17'd98830;
    value[878] = 17'd98828;
    value[879] = 17'd98825;
    value[880] = 17'd98822;
    value[881] = 17'd98820;
    value[882] = 17'd98817;
    value[883] = 17'd98814;
    value[884] = 17'd98812;
    value[885] = 17'd98809;
    value[886] = 17'd98806;
    value[887] = 17'd98804;
    value[888] = 17'd98801;
    value[889] = 17'd98798;
    value[890] = 17'd98795;
    value[891] = 17'd98793;
    value[892] = 17'd98790;
    value[893] = 17'd98787;
    value[894] = 17'd98785;
    value[895] = 17'd98782;
    value[896] = 17'd98779;
    value[897] = 17'd98777;
    value[898] = 17'd98774;
    value[899] = 17'd98771;
    value[900] = 17'd98768;
    value[901] = 17'd98766;
    value[902] = 17'd98763;
    value[903] = 17'd98760;
    value[904] = 17'd98757;
    value[905] = 17'd98755;
    value[906] = 17'd98752;
    value[907] = 17'd98749;
    value[908] = 17'd98746;
    value[909] = 17'd98744;
    value[910] = 17'd98741;
    value[911] = 17'd98738;
    value[912] = 17'd98735;
    value[913] = 17'd98733;
    value[914] = 17'd98730;
    value[915] = 17'd98727;
    value[916] = 17'd98724;
    value[917] = 17'd98721;
    value[918] = 17'd98719;
    value[919] = 17'd98716;
    value[920] = 17'd98713;
    value[921] = 17'd98710;
    value[922] = 17'd98708;
    value[923] = 17'd98705;
    value[924] = 17'd98702;
    value[925] = 17'd98699;
    value[926] = 17'd98696;
    value[927] = 17'd98694;
    value[928] = 17'd98691;
    value[929] = 17'd98688;
    value[930] = 17'd98685;
    value[931] = 17'd98682;
    value[932] = 17'd98679;
    value[933] = 17'd98677;
    value[934] = 17'd98674;
    value[935] = 17'd98671;
    value[936] = 17'd98668;
    value[937] = 17'd98665;
    value[938] = 17'd98662;
    value[939] = 17'd98660;
    value[940] = 17'd98657;
    value[941] = 17'd98654;
    value[942] = 17'd98651;
    value[943] = 17'd98648;
    value[944] = 17'd98645;
    value[945] = 17'd98642;
    value[946] = 17'd98640;
    value[947] = 17'd98637;
    value[948] = 17'd98634;
    value[949] = 17'd98631;
    value[950] = 17'd98628;
    value[951] = 17'd98625;
    value[952] = 17'd98622;
    value[953] = 17'd98619;
    value[954] = 17'd98617;
    value[955] = 17'd98614;
    value[956] = 17'd98611;
    value[957] = 17'd98608;
    value[958] = 17'd98605;
    value[959] = 17'd98602;
    value[960] = 17'd98599;
    value[961] = 17'd98596;
    value[962] = 17'd98593;
    value[963] = 17'd98590;
    value[964] = 17'd98587;
    value[965] = 17'd98585;
    value[966] = 17'd98582;
    value[967] = 17'd98579;
    value[968] = 17'd98576;
    value[969] = 17'd98573;
    value[970] = 17'd98570;
    value[971] = 17'd98567;
    value[972] = 17'd98564;
    value[973] = 17'd98561;
    value[974] = 17'd98558;
    value[975] = 17'd98555;
    value[976] = 17'd98552;
    value[977] = 17'd98549;
    value[978] = 17'd98546;
    value[979] = 17'd98543;
    value[980] = 17'd98540;
    value[981] = 17'd98537;
    value[982] = 17'd98534;
    value[983] = 17'd98531;
    value[984] = 17'd98528;
    value[985] = 17'd98525;
    value[986] = 17'd98522;
    value[987] = 17'd98519;
    value[988] = 17'd98516;
    value[989] = 17'd98513;
    value[990] = 17'd98510;
    value[991] = 17'd98507;
    value[992] = 17'd98504;
    value[993] = 17'd98501;
    value[994] = 17'd98498;
    value[995] = 17'd98495;
    value[996] = 17'd98492;
    value[997] = 17'd98489;
    value[998] = 17'd98486;
    value[999] = 17'd98483;
    value[1000] = 17'd98480;
    value[1001] = 17'd98477;
    value[1002] = 17'd98474;
    value[1003] = 17'd98471;
    value[1004] = 17'd98468;
    value[1005] = 17'd98465;
    value[1006] = 17'd98462;
    value[1007] = 17'd98459;
    value[1008] = 17'd98456;
    value[1009] = 17'd98453;
    value[1010] = 17'd98450;
    value[1011] = 17'd98447;
    value[1012] = 17'd98444;
    value[1013] = 17'd98441;
    value[1014] = 17'd98438;
    value[1015] = 17'd98434;
    value[1016] = 17'd98431;
    value[1017] = 17'd98428;
    value[1018] = 17'd98425;
    value[1019] = 17'd98422;
    value[1020] = 17'd98419;
    value[1021] = 17'd98416;
    value[1022] = 17'd98413;
    value[1023] = 17'd98410;
    value[1024] = 17'd98407;
    value[1025] = 17'd98404;
    value[1026] = 17'd98400;
    value[1027] = 17'd98397;
    value[1028] = 17'd98394;
    value[1029] = 17'd98391;
    value[1030] = 17'd98388;
    value[1031] = 17'd98385;
    value[1032] = 17'd98382;
    value[1033] = 17'd98379;
    value[1034] = 17'd98376;
    value[1035] = 17'd98372;
    value[1036] = 17'd98369;
    value[1037] = 17'd98366;
    value[1038] = 17'd98363;
    value[1039] = 17'd98360;
    value[1040] = 17'd98357;
    value[1041] = 17'd98353;
    value[1042] = 17'd98350;
    value[1043] = 17'd98347;
    value[1044] = 17'd98344;
    value[1045] = 17'd98341;
    value[1046] = 17'd98338;
    value[1047] = 17'd98335;
    value[1048] = 17'd98331;
    value[1049] = 17'd98328;
    value[1050] = 17'd98325;
    value[1051] = 17'd98322;
    value[1052] = 17'd98319;
    value[1053] = 17'd98315;
    value[1054] = 17'd98312;
    value[1055] = 17'd98309;
    value[1056] = 17'd98306;
    value[1057] = 17'd98303;
    value[1058] = 17'd98299;
    value[1059] = 17'd98296;
    value[1060] = 17'd98293;
    value[1061] = 17'd98290;
    value[1062] = 17'd98287;
    value[1063] = 17'd98283;
    value[1064] = 17'd98280;
    value[1065] = 17'd98277;
    value[1066] = 17'd98274;
    value[1067] = 17'd98270;
    value[1068] = 17'd98267;
    value[1069] = 17'd98264;
    value[1070] = 17'd98261;
    value[1071] = 17'd98258;
    value[1072] = 17'd98254;
    value[1073] = 17'd98251;
    value[1074] = 17'd98248;
    value[1075] = 17'd98245;
    value[1076] = 17'd98241;
    value[1077] = 17'd98238;
    value[1078] = 17'd98235;
    value[1079] = 17'd98231;
    value[1080] = 17'd98228;
    value[1081] = 17'd98225;
    value[1082] = 17'd98222;
    value[1083] = 17'd98218;
    value[1084] = 17'd98215;
    value[1085] = 17'd98212;
    value[1086] = 17'd98209;
    value[1087] = 17'd98205;
    value[1088] = 17'd98202;
    value[1089] = 17'd98199;
    value[1090] = 17'd98195;
    value[1091] = 17'd98192;
    value[1092] = 17'd98189;
    value[1093] = 17'd98185;
    value[1094] = 17'd98182;
    value[1095] = 17'd98179;
    value[1096] = 17'd98176;
    value[1097] = 17'd98172;
    value[1098] = 17'd98169;
    value[1099] = 17'd98166;
    value[1100] = 17'd98162;
    value[1101] = 17'd98159;
    value[1102] = 17'd98156;
    value[1103] = 17'd98152;
    value[1104] = 17'd98149;
    value[1105] = 17'd98146;
    value[1106] = 17'd98142;
    value[1107] = 17'd98139;
    value[1108] = 17'd98135;
    value[1109] = 17'd98132;
    value[1110] = 17'd98129;
    value[1111] = 17'd98125;
    value[1112] = 17'd98122;
    value[1113] = 17'd98119;
    value[1114] = 17'd98115;
    value[1115] = 17'd98112;
    value[1116] = 17'd98109;
    value[1117] = 17'd98105;
    value[1118] = 17'd98102;
    value[1119] = 17'd98098;
    value[1120] = 17'd98095;
    value[1121] = 17'd98092;
    value[1122] = 17'd98088;
    value[1123] = 17'd98085;
    value[1124] = 17'd98081;
    value[1125] = 17'd98078;
    value[1126] = 17'd98075;
    value[1127] = 17'd98071;
    value[1128] = 17'd98068;
    value[1129] = 17'd98064;
    value[1130] = 17'd98061;
    value[1131] = 17'd98058;
    value[1132] = 17'd98054;
    value[1133] = 17'd98051;
    value[1134] = 17'd98047;
    value[1135] = 17'd98044;
    value[1136] = 17'd98040;
    value[1137] = 17'd98037;
    value[1138] = 17'd98034;
    value[1139] = 17'd98030;
    value[1140] = 17'd98027;
    value[1141] = 17'd98023;
    value[1142] = 17'd98020;
    value[1143] = 17'd98016;
    value[1144] = 17'd98013;
    value[1145] = 17'd98009;
    value[1146] = 17'd98006;
    value[1147] = 17'd98002;
    value[1148] = 17'd97999;
    value[1149] = 17'd97995;
    value[1150] = 17'd97992;
    value[1151] = 17'd97988;
    value[1152] = 17'd97985;
    value[1153] = 17'd97982;
    value[1154] = 17'd97978;
    value[1155] = 17'd97975;
    value[1156] = 17'd97971;
    value[1157] = 17'd97968;
    value[1158] = 17'd97964;
    value[1159] = 17'd97961;
    value[1160] = 17'd97957;
    value[1161] = 17'd97954;
    value[1162] = 17'd97950;
    value[1163] = 17'd97946;
    value[1164] = 17'd97943;
    value[1165] = 17'd97939;
    value[1166] = 17'd97936;
    value[1167] = 17'd97932;
    value[1168] = 17'd97929;
    value[1169] = 17'd97925;
    value[1170] = 17'd97922;
    value[1171] = 17'd97918;
    value[1172] = 17'd97915;
    value[1173] = 17'd97911;
    value[1174] = 17'd97908;
    value[1175] = 17'd97904;
    value[1176] = 17'd97900;
    value[1177] = 17'd97897;
    value[1178] = 17'd97893;
    value[1179] = 17'd97890;
    value[1180] = 17'd97886;
    value[1181] = 17'd97883;
    value[1182] = 17'd97879;
    value[1183] = 17'd97876;
    value[1184] = 17'd97872;
    value[1185] = 17'd97868;
    value[1186] = 17'd97865;
    value[1187] = 17'd97861;
    value[1188] = 17'd97858;
    value[1189] = 17'd97854;
    value[1190] = 17'd97850;
    value[1191] = 17'd97847;
    value[1192] = 17'd97843;
    value[1193] = 17'd97840;
    value[1194] = 17'd97836;
    value[1195] = 17'd97832;
    value[1196] = 17'd97829;
    value[1197] = 17'd97825;
    value[1198] = 17'd97822;
    value[1199] = 17'd97818;
    value[1200] = 17'd97814;
    value[1201] = 17'd97811;
    value[1202] = 17'd97807;
    value[1203] = 17'd97803;
    value[1204] = 17'd97800;
    value[1205] = 17'd97796;
    value[1206] = 17'd97792;
    value[1207] = 17'd97789;
    value[1208] = 17'd97785;
    value[1209] = 17'd97781;
    value[1210] = 17'd97778;
    value[1211] = 17'd97774;
    value[1212] = 17'd97771;
    value[1213] = 17'd97767;
    value[1214] = 17'd97763;
    value[1215] = 17'd97759;
    value[1216] = 17'd97756;
    value[1217] = 17'd97752;
    value[1218] = 17'd97748;
    value[1219] = 17'd97745;
    value[1220] = 17'd97741;
    value[1221] = 17'd97737;
    value[1222] = 17'd97734;
    value[1223] = 17'd97730;
    value[1224] = 17'd97726;
    value[1225] = 17'd97723;
    value[1226] = 17'd97719;
    value[1227] = 17'd97715;
    value[1228] = 17'd97711;
    value[1229] = 17'd97708;
    value[1230] = 17'd97704;
    value[1231] = 17'd97700;
    value[1232] = 17'd97697;
    value[1233] = 17'd97693;
    value[1234] = 17'd97689;
    value[1235] = 17'd97685;
    value[1236] = 17'd97682;
    value[1237] = 17'd97678;
    value[1238] = 17'd97674;
    value[1239] = 17'd97670;
    value[1240] = 17'd97667;
    value[1241] = 17'd97663;
    value[1242] = 17'd97659;
    value[1243] = 17'd97655;
    value[1244] = 17'd97652;
    value[1245] = 17'd97648;
    value[1246] = 17'd97644;
    value[1247] = 17'd97640;
    value[1248] = 17'd97637;
    value[1249] = 17'd97633;
    value[1250] = 17'd97629;
    value[1251] = 17'd97625;
    value[1252] = 17'd97622;
    value[1253] = 17'd97618;
    value[1254] = 17'd97614;
    value[1255] = 17'd97610;
    value[1256] = 17'd97606;
    value[1257] = 17'd97603;
    value[1258] = 17'd97599;
    value[1259] = 17'd97595;
    value[1260] = 17'd97591;
    value[1261] = 17'd97587;
    value[1262] = 17'd97584;
    value[1263] = 17'd97580;
    value[1264] = 17'd97576;
    value[1265] = 17'd97572;
    value[1266] = 17'd97568;
    value[1267] = 17'd97564;
    value[1268] = 17'd97561;
    value[1269] = 17'd97557;
    value[1270] = 17'd97553;
    value[1271] = 17'd97549;
    value[1272] = 17'd97545;
    value[1273] = 17'd97541;
    value[1274] = 17'd97538;
    value[1275] = 17'd97534;
    value[1276] = 17'd97530;
    value[1277] = 17'd97526;
    value[1278] = 17'd97522;
    value[1279] = 17'd97518;
    value[1280] = 17'd97514;
    value[1281] = 17'd97511;
    value[1282] = 17'd97507;
    value[1283] = 17'd97503;
    value[1284] = 17'd97499;
    value[1285] = 17'd97495;
    value[1286] = 17'd97491;
    value[1287] = 17'd97487;
    value[1288] = 17'd97483;
    value[1289] = 17'd97480;
    value[1290] = 17'd97476;
    value[1291] = 17'd97472;
    value[1292] = 17'd97468;
    value[1293] = 17'd97464;
    value[1294] = 17'd97460;
    value[1295] = 17'd97456;
    value[1296] = 17'd97452;
    value[1297] = 17'd97448;
    value[1298] = 17'd97444;
    value[1299] = 17'd97440;
    value[1300] = 17'd97437;
    value[1301] = 17'd97433;
    value[1302] = 17'd97429;
    value[1303] = 17'd97425;
    value[1304] = 17'd97421;
    value[1305] = 17'd97417;
    value[1306] = 17'd97413;
    value[1307] = 17'd97409;
    value[1308] = 17'd97405;
    value[1309] = 17'd97401;
    value[1310] = 17'd97397;
    value[1311] = 17'd97393;
    value[1312] = 17'd97389;
    value[1313] = 17'd97385;
    value[1314] = 17'd97381;
    value[1315] = 17'd97377;
    value[1316] = 17'd97373;
    value[1317] = 17'd97369;
    value[1318] = 17'd97365;
    value[1319] = 17'd97361;
    value[1320] = 17'd97357;
    value[1321] = 17'd97353;
    value[1322] = 17'd97349;
    value[1323] = 17'd97345;
    value[1324] = 17'd97341;
    value[1325] = 17'd97337;
    value[1326] = 17'd97333;
    value[1327] = 17'd97329;
    value[1328] = 17'd97325;
    value[1329] = 17'd97321;
    value[1330] = 17'd97317;
    value[1331] = 17'd97313;
    value[1332] = 17'd97309;
    value[1333] = 17'd97305;
    value[1334] = 17'd97301;
    value[1335] = 17'd97297;
    value[1336] = 17'd97293;
    value[1337] = 17'd97289;
    value[1338] = 17'd97285;
    value[1339] = 17'd97281;
    value[1340] = 17'd97277;
    value[1341] = 17'd97273;
    value[1342] = 17'd97269;
    value[1343] = 17'd97265;
    value[1344] = 17'd97261;
    value[1345] = 17'd97257;
    value[1346] = 17'd97253;
    value[1347] = 17'd97249;
    value[1348] = 17'd97245;
    value[1349] = 17'd97241;
    value[1350] = 17'd97236;
    value[1351] = 17'd97232;
    value[1352] = 17'd97228;
    value[1353] = 17'd97224;
    value[1354] = 17'd97220;
    value[1355] = 17'd97216;
    value[1356] = 17'd97212;
    value[1357] = 17'd97208;
    value[1358] = 17'd97204;
    value[1359] = 17'd97200;
    value[1360] = 17'd97196;
    value[1361] = 17'd97191;
    value[1362] = 17'd97187;
    value[1363] = 17'd97183;
    value[1364] = 17'd97179;
    value[1365] = 17'd97175;
    value[1366] = 17'd97171;
    value[1367] = 17'd97167;
    value[1368] = 17'd97163;
    value[1369] = 17'd97159;
    value[1370] = 17'd97154;
    value[1371] = 17'd97150;
    value[1372] = 17'd97146;
    value[1373] = 17'd97142;
    value[1374] = 17'd97138;
    value[1375] = 17'd97134;
    value[1376] = 17'd97130;
    value[1377] = 17'd97125;
    value[1378] = 17'd97121;
    value[1379] = 17'd97117;
    value[1380] = 17'd97113;
    value[1381] = 17'd97109;
    value[1382] = 17'd97105;
    value[1383] = 17'd97100;
    value[1384] = 17'd97096;
    value[1385] = 17'd97092;
    value[1386] = 17'd97088;
    value[1387] = 17'd97084;
    value[1388] = 17'd97080;
    value[1389] = 17'd97075;
    value[1390] = 17'd97071;
    value[1391] = 17'd97067;
    value[1392] = 17'd97063;
    value[1393] = 17'd97059;
    value[1394] = 17'd97054;
    value[1395] = 17'd97050;
    value[1396] = 17'd97046;
    value[1397] = 17'd97042;
    value[1398] = 17'd97038;
    value[1399] = 17'd97033;
    value[1400] = 17'd97029;
    value[1401] = 17'd97025;
    value[1402] = 17'd97021;
    value[1403] = 17'd97016;
    value[1404] = 17'd97012;
    value[1405] = 17'd97008;
    value[1406] = 17'd97004;
    value[1407] = 17'd96999;
    value[1408] = 17'd96995;
    value[1409] = 17'd96991;
    value[1410] = 17'd96987;
    value[1411] = 17'd96982;
    value[1412] = 17'd96978;
    value[1413] = 17'd96974;
    value[1414] = 17'd96970;
    value[1415] = 17'd96965;
    value[1416] = 17'd96961;
    value[1417] = 17'd96957;
    value[1418] = 17'd96953;
    value[1419] = 17'd96948;
    value[1420] = 17'd96944;
    value[1421] = 17'd96940;
    value[1422] = 17'd96935;
    value[1423] = 17'd96931;
    value[1424] = 17'd96927;
    value[1425] = 17'd96923;
    value[1426] = 17'd96918;
    value[1427] = 17'd96914;
    value[1428] = 17'd96910;
    value[1429] = 17'd96905;
    value[1430] = 17'd96901;
    value[1431] = 17'd96897;
    value[1432] = 17'd96892;
    value[1433] = 17'd96888;
    value[1434] = 17'd96884;
    value[1435] = 17'd96879;
    value[1436] = 17'd96875;
    value[1437] = 17'd96871;
    value[1438] = 17'd96866;
    value[1439] = 17'd96862;
    value[1440] = 17'd96858;
    value[1441] = 17'd96853;
    value[1442] = 17'd96849;
    value[1443] = 17'd96845;
    value[1444] = 17'd96840;
    value[1445] = 17'd96836;
    value[1446] = 17'd96832;
    value[1447] = 17'd96827;
    value[1448] = 17'd96823;
    value[1449] = 17'd96819;
    value[1450] = 17'd96814;
    value[1451] = 17'd96810;
    value[1452] = 17'd96806;
    value[1453] = 17'd96801;
    value[1454] = 17'd96797;
    value[1455] = 17'd96792;
    value[1456] = 17'd96788;
    value[1457] = 17'd96784;
    value[1458] = 17'd96779;
    value[1459] = 17'd96775;
    value[1460] = 17'd96770;
    value[1461] = 17'd96766;
    value[1462] = 17'd96762;
    value[1463] = 17'd96757;
    value[1464] = 17'd96753;
    value[1465] = 17'd96748;
    value[1466] = 17'd96744;
    value[1467] = 17'd96740;
    value[1468] = 17'd96735;
    value[1469] = 17'd96731;
    value[1470] = 17'd96726;
    value[1471] = 17'd96722;
    value[1472] = 17'd96717;
    value[1473] = 17'd96713;
    value[1474] = 17'd96709;
    value[1475] = 17'd96704;
    value[1476] = 17'd96700;
    value[1477] = 17'd96695;
    value[1478] = 17'd96691;
    value[1479] = 17'd96686;
    value[1480] = 17'd96682;
    value[1481] = 17'd96677;
    value[1482] = 17'd96673;
    value[1483] = 17'd96668;
    value[1484] = 17'd96664;
    value[1485] = 17'd96660;
    value[1486] = 17'd96655;
    value[1487] = 17'd96651;
    value[1488] = 17'd96646;
    value[1489] = 17'd96642;
    value[1490] = 17'd96637;
    value[1491] = 17'd96633;
    value[1492] = 17'd96628;
    value[1493] = 17'd96624;
    value[1494] = 17'd96619;
    value[1495] = 17'd96615;
    value[1496] = 17'd96610;
    value[1497] = 17'd96606;
    value[1498] = 17'd96601;
    value[1499] = 17'd96597;
    value[1500] = 17'd96592;
    value[1501] = 17'd96588;
    value[1502] = 17'd96583;
    value[1503] = 17'd96579;
    value[1504] = 17'd96574;
    value[1505] = 17'd96569;
    value[1506] = 17'd96565;
    value[1507] = 17'd96560;
    value[1508] = 17'd96556;
    value[1509] = 17'd96551;
    value[1510] = 17'd96547;
    value[1511] = 17'd96542;
    value[1512] = 17'd96538;
    value[1513] = 17'd96533;
    value[1514] = 17'd96529;
    value[1515] = 17'd96524;
    value[1516] = 17'd96519;
    value[1517] = 17'd96515;
    value[1518] = 17'd96510;
    value[1519] = 17'd96506;
    value[1520] = 17'd96501;
    value[1521] = 17'd96497;
    value[1522] = 17'd96492;
    value[1523] = 17'd96487;
    value[1524] = 17'd96483;
    value[1525] = 17'd96478;
    value[1526] = 17'd96474;
    value[1527] = 17'd96469;
    value[1528] = 17'd96464;
    value[1529] = 17'd96460;
    value[1530] = 17'd96455;
    value[1531] = 17'd96451;
    value[1532] = 17'd96446;
    value[1533] = 17'd96441;
    value[1534] = 17'd96437;
    value[1535] = 17'd96432;
    value[1536] = 17'd96428;
    value[1537] = 17'd96423;
    value[1538] = 17'd96418;
    value[1539] = 17'd96414;
    value[1540] = 17'd96409;
    value[1541] = 17'd96404;
    value[1542] = 17'd96400;
    value[1543] = 17'd96395;
    value[1544] = 17'd96390;
    value[1545] = 17'd96386;
    value[1546] = 17'd96381;
    value[1547] = 17'd96377;
    value[1548] = 17'd96372;
    value[1549] = 17'd96367;
    value[1550] = 17'd96363;
    value[1551] = 17'd96358;
    value[1552] = 17'd96353;
    value[1553] = 17'd96349;
    value[1554] = 17'd96344;
    value[1555] = 17'd96339;
    value[1556] = 17'd96335;
    value[1557] = 17'd96330;
    value[1558] = 17'd96325;
    value[1559] = 17'd96320;
    value[1560] = 17'd96316;
    value[1561] = 17'd96311;
    value[1562] = 17'd96306;
    value[1563] = 17'd96302;
    value[1564] = 17'd96297;
    value[1565] = 17'd96292;
    value[1566] = 17'd96288;
    value[1567] = 17'd96283;
    value[1568] = 17'd96278;
    value[1569] = 17'd96273;
    value[1570] = 17'd96269;
    value[1571] = 17'd96264;
    value[1572] = 17'd96259;
    value[1573] = 17'd96254;
    value[1574] = 17'd96250;
    value[1575] = 17'd96245;
    value[1576] = 17'd96240;
    value[1577] = 17'd96236;
    value[1578] = 17'd96231;
    value[1579] = 17'd96226;
    value[1580] = 17'd96221;
    value[1581] = 17'd96217;
    value[1582] = 17'd96212;
    value[1583] = 17'd96207;
    value[1584] = 17'd96202;
    value[1585] = 17'd96198;
    value[1586] = 17'd96193;
    value[1587] = 17'd96188;
    value[1588] = 17'd96183;
    value[1589] = 17'd96178;
    value[1590] = 17'd96174;
    value[1591] = 17'd96169;
    value[1592] = 17'd96164;
    value[1593] = 17'd96159;
    value[1594] = 17'd96154;
    value[1595] = 17'd96150;
    value[1596] = 17'd96145;
    value[1597] = 17'd96140;
    value[1598] = 17'd96135;
    value[1599] = 17'd96130;
    value[1600] = 17'd96126;
    value[1601] = 17'd96121;
    value[1602] = 17'd96116;
    value[1603] = 17'd96111;
    value[1604] = 17'd96106;
    value[1605] = 17'd96102;
    value[1606] = 17'd96097;
    value[1607] = 17'd96092;
    value[1608] = 17'd96087;
    value[1609] = 17'd96082;
    value[1610] = 17'd96077;
    value[1611] = 17'd96073;
    value[1612] = 17'd96068;
    value[1613] = 17'd96063;
    value[1614] = 17'd96058;
    value[1615] = 17'd96053;
    value[1616] = 17'd96048;
    value[1617] = 17'd96043;
    value[1618] = 17'd96039;
    value[1619] = 17'd96034;
    value[1620] = 17'd96029;
    value[1621] = 17'd96024;
    value[1622] = 17'd96019;
    value[1623] = 17'd96014;
    value[1624] = 17'd96009;
    value[1625] = 17'd96004;
    value[1626] = 17'd96000;
    value[1627] = 17'd95995;
    value[1628] = 17'd95990;
    value[1629] = 17'd95985;
    value[1630] = 17'd95980;
    value[1631] = 17'd95975;
    value[1632] = 17'd95970;
    value[1633] = 17'd95965;
    value[1634] = 17'd95960;
    value[1635] = 17'd95956;
    value[1636] = 17'd95951;
    value[1637] = 17'd95946;
    value[1638] = 17'd95941;
    value[1639] = 17'd95936;
    value[1640] = 17'd95931;
    value[1641] = 17'd95926;
    value[1642] = 17'd95921;
    value[1643] = 17'd95916;
    value[1644] = 17'd95911;
    value[1645] = 17'd95906;
    value[1646] = 17'd95901;
    value[1647] = 17'd95896;
    value[1648] = 17'd95891;
    value[1649] = 17'd95886;
    value[1650] = 17'd95881;
    value[1651] = 17'd95877;
    value[1652] = 17'd95872;
    value[1653] = 17'd95867;
    value[1654] = 17'd95862;
    value[1655] = 17'd95857;
    value[1656] = 17'd95852;
    value[1657] = 17'd95847;
    value[1658] = 17'd95842;
    value[1659] = 17'd95837;
    value[1660] = 17'd95832;
    value[1661] = 17'd95827;
    value[1662] = 17'd95822;
    value[1663] = 17'd95817;
    value[1664] = 17'd95812;
    value[1665] = 17'd95807;
    value[1666] = 17'd95802;
    value[1667] = 17'd95797;
    value[1668] = 17'd95792;
    value[1669] = 17'd95787;
    value[1670] = 17'd95782;
    value[1671] = 17'd95777;
    value[1672] = 17'd95772;
    value[1673] = 17'd95767;
    value[1674] = 17'd95762;
    value[1675] = 17'd95757;
    value[1676] = 17'd95752;
    value[1677] = 17'd95747;
    value[1678] = 17'd95742;
    value[1679] = 17'd95736;
    value[1680] = 17'd95731;
    value[1681] = 17'd95726;
    value[1682] = 17'd95721;
    value[1683] = 17'd95716;
    value[1684] = 17'd95711;
    value[1685] = 17'd95706;
    value[1686] = 17'd95701;
    value[1687] = 17'd95696;
    value[1688] = 17'd95691;
    value[1689] = 17'd95686;
    value[1690] = 17'd95681;
    value[1691] = 17'd95676;
    value[1692] = 17'd95671;
    value[1693] = 17'd95666;
    value[1694] = 17'd95661;
    value[1695] = 17'd95655;
    value[1696] = 17'd95650;
    value[1697] = 17'd95645;
    value[1698] = 17'd95640;
    value[1699] = 17'd95635;
    value[1700] = 17'd95630;
    value[1701] = 17'd95625;
    value[1702] = 17'd95620;
    value[1703] = 17'd95615;
    value[1704] = 17'd95610;
    value[1705] = 17'd95604;
    value[1706] = 17'd95599;
    value[1707] = 17'd95594;
    value[1708] = 17'd95589;
    value[1709] = 17'd95584;
    value[1710] = 17'd95579;
    value[1711] = 17'd95574;
    value[1712] = 17'd95569;
    value[1713] = 17'd95563;
    value[1714] = 17'd95558;
    value[1715] = 17'd95553;
    value[1716] = 17'd95548;
    value[1717] = 17'd95543;
    value[1718] = 17'd95538;
    value[1719] = 17'd95532;
    value[1720] = 17'd95527;
    value[1721] = 17'd95522;
    value[1722] = 17'd95517;
    value[1723] = 17'd95512;
    value[1724] = 17'd95507;
    value[1725] = 17'd95501;
    value[1726] = 17'd95496;
    value[1727] = 17'd95491;
    value[1728] = 17'd95486;
    value[1729] = 17'd95481;
    value[1730] = 17'd95476;
    value[1731] = 17'd95470;
    value[1732] = 17'd95465;
    value[1733] = 17'd95460;
    value[1734] = 17'd95455;
    value[1735] = 17'd95450;
    value[1736] = 17'd95444;
    value[1737] = 17'd95439;
    value[1738] = 17'd95434;
    value[1739] = 17'd95429;
    value[1740] = 17'd95424;
    value[1741] = 17'd95418;
    value[1742] = 17'd95413;
    value[1743] = 17'd95408;
    value[1744] = 17'd95403;
    value[1745] = 17'd95397;
    value[1746] = 17'd95392;
    value[1747] = 17'd95387;
    value[1748] = 17'd95382;
    value[1749] = 17'd95376;
    value[1750] = 17'd95371;
    value[1751] = 17'd95366;
    value[1752] = 17'd95361;
    value[1753] = 17'd95355;
    value[1754] = 17'd95350;
    value[1755] = 17'd95345;
    value[1756] = 17'd95340;
    value[1757] = 17'd95334;
    value[1758] = 17'd95329;
    value[1759] = 17'd95324;
    value[1760] = 17'd95319;
    value[1761] = 17'd95313;
    value[1762] = 17'd95308;
    value[1763] = 17'd95303;
    value[1764] = 17'd95297;
    value[1765] = 17'd95292;
    value[1766] = 17'd95287;
    value[1767] = 17'd95282;
    value[1768] = 17'd95276;
    value[1769] = 17'd95271;
    value[1770] = 17'd95266;
    value[1771] = 17'd95260;
    value[1772] = 17'd95255;
    value[1773] = 17'd95250;
    value[1774] = 17'd95244;
    value[1775] = 17'd95239;
    value[1776] = 17'd95234;
    value[1777] = 17'd95228;
    value[1778] = 17'd95223;
    value[1779] = 17'd95218;
    value[1780] = 17'd95212;
    value[1781] = 17'd95207;
    value[1782] = 17'd95202;
    value[1783] = 17'd95196;
    value[1784] = 17'd95191;
    value[1785] = 17'd95186;
    value[1786] = 17'd95180;
    value[1787] = 17'd95175;
    value[1788] = 17'd95170;
    value[1789] = 17'd95164;
    value[1790] = 17'd95159;
    value[1791] = 17'd95154;
    value[1792] = 17'd95148;
    value[1793] = 17'd95143;
    value[1794] = 17'd95137;
    value[1795] = 17'd95132;
    value[1796] = 17'd95127;
    value[1797] = 17'd95121;
    value[1798] = 17'd95116;
    value[1799] = 17'd95111;
    value[1800] = 17'd95105;
    value[1801] = 17'd95100;
    value[1802] = 17'd95094;
    value[1803] = 17'd95089;
    value[1804] = 17'd95084;
    value[1805] = 17'd95078;
    value[1806] = 17'd95073;
    value[1807] = 17'd95067;
    value[1808] = 17'd95062;
    value[1809] = 17'd95056;
    value[1810] = 17'd95051;
    value[1811] = 17'd95046;
    value[1812] = 17'd95040;
    value[1813] = 17'd95035;
    value[1814] = 17'd95029;
    value[1815] = 17'd95024;
    value[1816] = 17'd95018;
    value[1817] = 17'd95013;
    value[1818] = 17'd95008;
    value[1819] = 17'd95002;
    value[1820] = 17'd94997;
    value[1821] = 17'd94991;
    value[1822] = 17'd94986;
    value[1823] = 17'd94980;
    value[1824] = 17'd94975;
    value[1825] = 17'd94969;
    value[1826] = 17'd94964;
    value[1827] = 17'd94958;
    value[1828] = 17'd94953;
    value[1829] = 17'd94948;
    value[1830] = 17'd94942;
    value[1831] = 17'd94937;
    value[1832] = 17'd94931;
    value[1833] = 17'd94926;
    value[1834] = 17'd94920;
    value[1835] = 17'd94915;
    value[1836] = 17'd94909;
    value[1837] = 17'd94904;
    value[1838] = 17'd94898;
    value[1839] = 17'd94893;
    value[1840] = 17'd94887;
    value[1841] = 17'd94882;
    value[1842] = 17'd94876;
    value[1843] = 17'd94871;
    value[1844] = 17'd94865;
    value[1845] = 17'd94860;
    value[1846] = 17'd94854;
    value[1847] = 17'd94848;
    value[1848] = 17'd94843;
    value[1849] = 17'd94837;
    value[1850] = 17'd94832;
    value[1851] = 17'd94826;
    value[1852] = 17'd94821;
    value[1853] = 17'd94815;
    value[1854] = 17'd94810;
    value[1855] = 17'd94804;
    value[1856] = 17'd94799;
    value[1857] = 17'd94793;
    value[1858] = 17'd94787;
    value[1859] = 17'd94782;
    value[1860] = 17'd94776;
    value[1861] = 17'd94771;
    value[1862] = 17'd94765;
    value[1863] = 17'd94760;
    value[1864] = 17'd94754;
    value[1865] = 17'd94748;
    value[1866] = 17'd94743;
    value[1867] = 17'd94737;
    value[1868] = 17'd94732;
    value[1869] = 17'd94726;
    value[1870] = 17'd94721;
    value[1871] = 17'd94715;
    value[1872] = 17'd94709;
    value[1873] = 17'd94704;
    value[1874] = 17'd94698;
    value[1875] = 17'd94693;
    value[1876] = 17'd94687;
    value[1877] = 17'd94681;
    value[1878] = 17'd94676;
    value[1879] = 17'd94670;
    value[1880] = 17'd94664;
    value[1881] = 17'd94659;
    value[1882] = 17'd94653;
    value[1883] = 17'd94648;
    value[1884] = 17'd94642;
    value[1885] = 17'd94636;
    value[1886] = 17'd94631;
    value[1887] = 17'd94625;
    value[1888] = 17'd94619;
    value[1889] = 17'd94614;
    value[1890] = 17'd94608;
    value[1891] = 17'd94602;
    value[1892] = 17'd94597;
    value[1893] = 17'd94591;
    value[1894] = 17'd94585;
    value[1895] = 17'd94580;
    value[1896] = 17'd94574;
    value[1897] = 17'd94568;
    value[1898] = 17'd94563;
    value[1899] = 17'd94557;
    value[1900] = 17'd94551;
    value[1901] = 17'd94546;
    value[1902] = 17'd94540;
    value[1903] = 17'd94534;
    value[1904] = 17'd94529;
    value[1905] = 17'd94523;
    value[1906] = 17'd94517;
    value[1907] = 17'd94512;
    value[1908] = 17'd94506;
    value[1909] = 17'd94500;
    value[1910] = 17'd94494;
    value[1911] = 17'd94489;
    value[1912] = 17'd94483;
    value[1913] = 17'd94477;
    value[1914] = 17'd94472;
    value[1915] = 17'd94466;
    value[1916] = 17'd94460;
    value[1917] = 17'd94454;
    value[1918] = 17'd94449;
    value[1919] = 17'd94443;
    value[1920] = 17'd94437;
    value[1921] = 17'd94431;
    value[1922] = 17'd94426;
    value[1923] = 17'd94420;
    value[1924] = 17'd94414;
    value[1925] = 17'd94408;
    value[1926] = 17'd94403;
    value[1927] = 17'd94397;
    value[1928] = 17'd94391;
    value[1929] = 17'd94385;
    value[1930] = 17'd94380;
    value[1931] = 17'd94374;
    value[1932] = 17'd94368;
    value[1933] = 17'd94362;
    value[1934] = 17'd94357;
    value[1935] = 17'd94351;
    value[1936] = 17'd94345;
    value[1937] = 17'd94339;
    value[1938] = 17'd94333;
    value[1939] = 17'd94328;
    value[1940] = 17'd94322;
    value[1941] = 17'd94316;
    value[1942] = 17'd94310;
    value[1943] = 17'd94304;
    value[1944] = 17'd94299;
    value[1945] = 17'd94293;
    value[1946] = 17'd94287;
    value[1947] = 17'd94281;
    value[1948] = 17'd94275;
    value[1949] = 17'd94269;
    value[1950] = 17'd94264;
    value[1951] = 17'd94258;
    value[1952] = 17'd94252;
    value[1953] = 17'd94246;
    value[1954] = 17'd94240;
    value[1955] = 17'd94234;
    value[1956] = 17'd94229;
    value[1957] = 17'd94223;
    value[1958] = 17'd94217;
    value[1959] = 17'd94211;
    value[1960] = 17'd94205;
    value[1961] = 17'd94199;
    value[1962] = 17'd94194;
    value[1963] = 17'd94188;
    value[1964] = 17'd94182;
    value[1965] = 17'd94176;
    value[1966] = 17'd94170;
    value[1967] = 17'd94164;
    value[1968] = 17'd94158;
    value[1969] = 17'd94152;
    value[1970] = 17'd94147;
    value[1971] = 17'd94141;
    value[1972] = 17'd94135;
    value[1973] = 17'd94129;
    value[1974] = 17'd94123;
    value[1975] = 17'd94117;
    value[1976] = 17'd94111;
    value[1977] = 17'd94105;
    value[1978] = 17'd94099;
    value[1979] = 17'd94093;
    value[1980] = 17'd94088;
    value[1981] = 17'd94082;
    value[1982] = 17'd94076;
    value[1983] = 17'd94070;
    value[1984] = 17'd94064;
    value[1985] = 17'd94058;
    value[1986] = 17'd94052;
    value[1987] = 17'd94046;
    value[1988] = 17'd94040;
    value[1989] = 17'd94034;
    value[1990] = 17'd94028;
    value[1991] = 17'd94022;
    value[1992] = 17'd94016;
    value[1993] = 17'd94010;
    value[1994] = 17'd94005;
    value[1995] = 17'd93999;
    value[1996] = 17'd93993;
    value[1997] = 17'd93987;
    value[1998] = 17'd93981;
    value[1999] = 17'd93975;
    value[2000] = 17'd93969;
    value[2001] = 17'd93963;
    value[2002] = 17'd93957;
    value[2003] = 17'd93951;
    value[2004] = 17'd93945;
    value[2005] = 17'd93939;
    value[2006] = 17'd93933;
    value[2007] = 17'd93927;
    value[2008] = 17'd93921;
    value[2009] = 17'd93915;
    value[2010] = 17'd93909;
    value[2011] = 17'd93903;
    value[2012] = 17'd93897;
    value[2013] = 17'd93891;
    value[2014] = 17'd93885;
    value[2015] = 17'd93879;
    value[2016] = 17'd93873;
    value[2017] = 17'd93867;
    value[2018] = 17'd93861;
    value[2019] = 17'd93855;
    value[2020] = 17'd93849;
    value[2021] = 17'd93843;
    value[2022] = 17'd93837;
    value[2023] = 17'd93831;
    value[2024] = 17'd93825;
    value[2025] = 17'd93819;
    value[2026] = 17'd93813;
    value[2027] = 17'd93807;
    value[2028] = 17'd93801;
    value[2029] = 17'd93794;
    value[2030] = 17'd93788;
    value[2031] = 17'd93782;
    value[2032] = 17'd93776;
    value[2033] = 17'd93770;
    value[2034] = 17'd93764;
    value[2035] = 17'd93758;
    value[2036] = 17'd93752;
    value[2037] = 17'd93746;
    value[2038] = 17'd93740;
    value[2039] = 17'd93734;
    value[2040] = 17'd93728;
    value[2041] = 17'd93722;
    value[2042] = 17'd93716;
    value[2043] = 17'd93709;
    value[2044] = 17'd93703;
    value[2045] = 17'd93697;
    value[2046] = 17'd93691;
    value[2047] = 17'd93685;
    value[2048] = 17'd93679;
    value[2049] = 17'd93673;
    value[2050] = 17'd93667;
    value[2051] = 17'd93661;
    value[2052] = 17'd93654;
    value[2053] = 17'd93648;
    value[2054] = 17'd93642;
    value[2055] = 17'd93636;
    value[2056] = 17'd93630;
    value[2057] = 17'd93624;
    value[2058] = 17'd93618;
    value[2059] = 17'd93612;
    value[2060] = 17'd93605;
    value[2061] = 17'd93599;
    value[2062] = 17'd93593;
    value[2063] = 17'd93587;
    value[2064] = 17'd93581;
    value[2065] = 17'd93575;
    value[2066] = 17'd93569;
    value[2067] = 17'd93562;
    value[2068] = 17'd93556;
    value[2069] = 17'd93550;
    value[2070] = 17'd93544;
    value[2071] = 17'd93538;
    value[2072] = 17'd93532;
    value[2073] = 17'd93525;
    value[2074] = 17'd93519;
    value[2075] = 17'd93513;
    value[2076] = 17'd93507;
    value[2077] = 17'd93501;
    value[2078] = 17'd93494;
    value[2079] = 17'd93488;
    value[2080] = 17'd93482;
    value[2081] = 17'd93476;
    value[2082] = 17'd93470;
    value[2083] = 17'd93463;
    value[2084] = 17'd93457;
    value[2085] = 17'd93451;
    value[2086] = 17'd93445;
    value[2087] = 17'd93439;
    value[2088] = 17'd93432;
    value[2089] = 17'd93426;
    value[2090] = 17'd93420;
    value[2091] = 17'd93414;
    value[2092] = 17'd93407;
    value[2093] = 17'd93401;
    value[2094] = 17'd93395;
    value[2095] = 17'd93389;
    value[2096] = 17'd93383;
    value[2097] = 17'd93376;
    value[2098] = 17'd93370;
    value[2099] = 17'd93364;
    value[2100] = 17'd93358;
    value[2101] = 17'd93351;
    value[2102] = 17'd93345;
    value[2103] = 17'd93339;
    value[2104] = 17'd93333;
    value[2105] = 17'd93326;
    value[2106] = 17'd93320;
    value[2107] = 17'd93314;
    value[2108] = 17'd93307;
    value[2109] = 17'd93301;
    value[2110] = 17'd93295;
    value[2111] = 17'd93289;
    value[2112] = 17'd93282;
    value[2113] = 17'd93276;
    value[2114] = 17'd93270;
    value[2115] = 17'd93263;
    value[2116] = 17'd93257;
    value[2117] = 17'd93251;
    value[2118] = 17'd93245;
    value[2119] = 17'd93238;
    value[2120] = 17'd93232;
    value[2121] = 17'd93226;
    value[2122] = 17'd93219;
    value[2123] = 17'd93213;
    value[2124] = 17'd93207;
    value[2125] = 17'd93200;
    value[2126] = 17'd93194;
    value[2127] = 17'd93188;
    value[2128] = 17'd93181;
    value[2129] = 17'd93175;
    value[2130] = 17'd93169;
    value[2131] = 17'd93162;
    value[2132] = 17'd93156;
    value[2133] = 17'd93150;
    value[2134] = 17'd93143;
    value[2135] = 17'd93137;
    value[2136] = 17'd93131;
    value[2137] = 17'd93124;
    value[2138] = 17'd93118;
    value[2139] = 17'd93111;
    value[2140] = 17'd93105;
    value[2141] = 17'd93099;
    value[2142] = 17'd93092;
    value[2143] = 17'd93086;
    value[2144] = 17'd93080;
    value[2145] = 17'd93073;
    value[2146] = 17'd93067;
    value[2147] = 17'd93060;
    value[2148] = 17'd93054;
    value[2149] = 17'd93048;
    value[2150] = 17'd93041;
    value[2151] = 17'd93035;
    value[2152] = 17'd93028;
    value[2153] = 17'd93022;
    value[2154] = 17'd93016;
    value[2155] = 17'd93009;
    value[2156] = 17'd93003;
    value[2157] = 17'd92996;
    value[2158] = 17'd92990;
    value[2159] = 17'd92984;
    value[2160] = 17'd92977;
    value[2161] = 17'd92971;
    value[2162] = 17'd92964;
    value[2163] = 17'd92958;
    value[2164] = 17'd92951;
    value[2165] = 17'd92945;
    value[2166] = 17'd92939;
    value[2167] = 17'd92932;
    value[2168] = 17'd92926;
    value[2169] = 17'd92919;
    value[2170] = 17'd92913;
    value[2171] = 17'd92906;
    value[2172] = 17'd92900;
    value[2173] = 17'd92893;
    value[2174] = 17'd92887;
    value[2175] = 17'd92880;
    value[2176] = 17'd92874;
    value[2177] = 17'd92868;
    value[2178] = 17'd92861;
    value[2179] = 17'd92855;
    value[2180] = 17'd92848;
    value[2181] = 17'd92842;
    value[2182] = 17'd92835;
    value[2183] = 17'd92829;
    value[2184] = 17'd92822;
    value[2185] = 17'd92816;
    value[2186] = 17'd92809;
    value[2187] = 17'd92803;
    value[2188] = 17'd92796;
    value[2189] = 17'd92790;
    value[2190] = 17'd92783;
    value[2191] = 17'd92777;
    value[2192] = 17'd92770;
    value[2193] = 17'd92764;
    value[2194] = 17'd92757;
    value[2195] = 17'd92751;
    value[2196] = 17'd92744;
    value[2197] = 17'd92737;
    value[2198] = 17'd92731;
    value[2199] = 17'd92724;
    value[2200] = 17'd92718;
    value[2201] = 17'd92711;
    value[2202] = 17'd92705;
    value[2203] = 17'd92698;
    value[2204] = 17'd92692;
    value[2205] = 17'd92685;
    value[2206] = 17'd92679;
    value[2207] = 17'd92672;
    value[2208] = 17'd92665;
    value[2209] = 17'd92659;
    value[2210] = 17'd92652;
    value[2211] = 17'd92646;
    value[2212] = 17'd92639;
    value[2213] = 17'd92633;
    value[2214] = 17'd92626;
    value[2215] = 17'd92619;
    value[2216] = 17'd92613;
    value[2217] = 17'd92606;
    value[2218] = 17'd92600;
    value[2219] = 17'd92593;
    value[2220] = 17'd92587;
    value[2221] = 17'd92580;
    value[2222] = 17'd92573;
    value[2223] = 17'd92567;
    value[2224] = 17'd92560;
    value[2225] = 17'd92554;
    value[2226] = 17'd92547;
    value[2227] = 17'd92540;
    value[2228] = 17'd92534;
    value[2229] = 17'd92527;
    value[2230] = 17'd92520;
    value[2231] = 17'd92514;
    value[2232] = 17'd92507;
    value[2233] = 17'd92501;
    value[2234] = 17'd92494;
    value[2235] = 17'd92487;
    value[2236] = 17'd92481;
    value[2237] = 17'd92474;
    value[2238] = 17'd92467;
    value[2239] = 17'd92461;
    value[2240] = 17'd92454;
    value[2241] = 17'd92447;
    value[2242] = 17'd92441;
    value[2243] = 17'd92434;
    value[2244] = 17'd92427;
    value[2245] = 17'd92421;
    value[2246] = 17'd92414;
    value[2247] = 17'd92407;
    value[2248] = 17'd92401;
    value[2249] = 17'd92394;
    value[2250] = 17'd92387;
    value[2251] = 17'd92381;
    value[2252] = 17'd92374;
    value[2253] = 17'd92367;
    value[2254] = 17'd92361;
    value[2255] = 17'd92354;
    value[2256] = 17'd92347;
    value[2257] = 17'd92341;
    value[2258] = 17'd92334;
    value[2259] = 17'd92327;
    value[2260] = 17'd92321;
    value[2261] = 17'd92314;
    value[2262] = 17'd92307;
    value[2263] = 17'd92300;
    value[2264] = 17'd92294;
    value[2265] = 17'd92287;
    value[2266] = 17'd92280;
    value[2267] = 17'd92274;
    value[2268] = 17'd92267;
    value[2269] = 17'd92260;
    value[2270] = 17'd92253;
    value[2271] = 17'd92247;
    value[2272] = 17'd92240;
    value[2273] = 17'd92233;
    value[2274] = 17'd92226;
    value[2275] = 17'd92220;
    value[2276] = 17'd92213;
    value[2277] = 17'd92206;
    value[2278] = 17'd92199;
    value[2279] = 17'd92193;
    value[2280] = 17'd92186;
    value[2281] = 17'd92179;
    value[2282] = 17'd92172;
    value[2283] = 17'd92166;
    value[2284] = 17'd92159;
    value[2285] = 17'd92152;
    value[2286] = 17'd92145;
    value[2287] = 17'd92138;
    value[2288] = 17'd92132;
    value[2289] = 17'd92125;
    value[2290] = 17'd92118;
    value[2291] = 17'd92111;
    value[2292] = 17'd92104;
    value[2293] = 17'd92098;
    value[2294] = 17'd92091;
    value[2295] = 17'd92084;
    value[2296] = 17'd92077;
    value[2297] = 17'd92070;
    value[2298] = 17'd92064;
    value[2299] = 17'd92057;
    value[2300] = 17'd92050;
    value[2301] = 17'd92043;
    value[2302] = 17'd92036;
    value[2303] = 17'd92030;
    value[2304] = 17'd92023;
    value[2305] = 17'd92016;
    value[2306] = 17'd92009;
    value[2307] = 17'd92002;
    value[2308] = 17'd91995;
    value[2309] = 17'd91988;
    value[2310] = 17'd91982;
    value[2311] = 17'd91975;
    value[2312] = 17'd91968;
    value[2313] = 17'd91961;
    value[2314] = 17'd91954;
    value[2315] = 17'd91947;
    value[2316] = 17'd91941;
    value[2317] = 17'd91934;
    value[2318] = 17'd91927;
    value[2319] = 17'd91920;
    value[2320] = 17'd91913;
    value[2321] = 17'd91906;
    value[2322] = 17'd91899;
    value[2323] = 17'd91892;
    value[2324] = 17'd91886;
    value[2325] = 17'd91879;
    value[2326] = 17'd91872;
    value[2327] = 17'd91865;
    value[2328] = 17'd91858;
    value[2329] = 17'd91851;
    value[2330] = 17'd91844;
    value[2331] = 17'd91837;
    value[2332] = 17'd91830;
    value[2333] = 17'd91823;
    value[2334] = 17'd91817;
    value[2335] = 17'd91810;
    value[2336] = 17'd91803;
    value[2337] = 17'd91796;
    value[2338] = 17'd91789;
    value[2339] = 17'd91782;
    value[2340] = 17'd91775;
    value[2341] = 17'd91768;
    value[2342] = 17'd91761;
    value[2343] = 17'd91754;
    value[2344] = 17'd91747;
    value[2345] = 17'd91740;
    value[2346] = 17'd91733;
    value[2347] = 17'd91726;
    value[2348] = 17'd91719;
    value[2349] = 17'd91712;
    value[2350] = 17'd91706;
    value[2351] = 17'd91699;
    value[2352] = 17'd91692;
    value[2353] = 17'd91685;
    value[2354] = 17'd91678;
    value[2355] = 17'd91671;
    value[2356] = 17'd91664;
    value[2357] = 17'd91657;
    value[2358] = 17'd91650;
    value[2359] = 17'd91643;
    value[2360] = 17'd91636;
    value[2361] = 17'd91629;
    value[2362] = 17'd91622;
    value[2363] = 17'd91615;
    value[2364] = 17'd91608;
    value[2365] = 17'd91601;
    value[2366] = 17'd91594;
    value[2367] = 17'd91587;
    value[2368] = 17'd91580;
    value[2369] = 17'd91573;
    value[2370] = 17'd91566;
    value[2371] = 17'd91559;
    value[2372] = 17'd91552;
    value[2373] = 17'd91545;
    value[2374] = 17'd91538;
    value[2375] = 17'd91531;
    value[2376] = 17'd91524;
    value[2377] = 17'd91517;
    value[2378] = 17'd91510;
    value[2379] = 17'd91503;
    value[2380] = 17'd91495;
    value[2381] = 17'd91488;
    value[2382] = 17'd91481;
    value[2383] = 17'd91474;
    value[2384] = 17'd91467;
    value[2385] = 17'd91460;
    value[2386] = 17'd91453;
    value[2387] = 17'd91446;
    value[2388] = 17'd91439;
    value[2389] = 17'd91432;
    value[2390] = 17'd91425;
    value[2391] = 17'd91418;
    value[2392] = 17'd91411;
    value[2393] = 17'd91404;
    value[2394] = 17'd91397;
    value[2395] = 17'd91390;
    value[2396] = 17'd91382;
    value[2397] = 17'd91375;
    value[2398] = 17'd91368;
    value[2399] = 17'd91361;
    value[2400] = 17'd91354;
    value[2401] = 17'd91347;
    value[2402] = 17'd91340;
    value[2403] = 17'd91333;
    value[2404] = 17'd91326;
    value[2405] = 17'd91319;
    value[2406] = 17'd91311;
    value[2407] = 17'd91304;
    value[2408] = 17'd91297;
    value[2409] = 17'd91290;
    value[2410] = 17'd91283;
    value[2411] = 17'd91276;
    value[2412] = 17'd91269;
    value[2413] = 17'd91262;
    value[2414] = 17'd91254;
    value[2415] = 17'd91247;
    value[2416] = 17'd91240;
    value[2417] = 17'd91233;
    value[2418] = 17'd91226;
    value[2419] = 17'd91219;
    value[2420] = 17'd91212;
    value[2421] = 17'd91204;
    value[2422] = 17'd91197;
    value[2423] = 17'd91190;
    value[2424] = 17'd91183;
    value[2425] = 17'd91176;
    value[2426] = 17'd91169;
    value[2427] = 17'd91161;
    value[2428] = 17'd91154;
    value[2429] = 17'd91147;
    value[2430] = 17'd91140;
    value[2431] = 17'd91133;
    value[2432] = 17'd91125;
    value[2433] = 17'd91118;
    value[2434] = 17'd91111;
    value[2435] = 17'd91104;
    value[2436] = 17'd91097;
    value[2437] = 17'd91089;
    value[2438] = 17'd91082;
    value[2439] = 17'd91075;
    value[2440] = 17'd91068;
    value[2441] = 17'd91061;
    value[2442] = 17'd91053;
    value[2443] = 17'd91046;
    value[2444] = 17'd91039;
    value[2445] = 17'd91032;
    value[2446] = 17'd91025;
    value[2447] = 17'd91017;
    value[2448] = 17'd91010;
    value[2449] = 17'd91003;
    value[2450] = 17'd90996;
    value[2451] = 17'd90988;
    value[2452] = 17'd90981;
    value[2453] = 17'd90974;
    value[2454] = 17'd90967;
    value[2455] = 17'd90959;
    value[2456] = 17'd90952;
    value[2457] = 17'd90945;
    value[2458] = 17'd90938;
    value[2459] = 17'd90930;
    value[2460] = 17'd90923;
    value[2461] = 17'd90916;
    value[2462] = 17'd90909;
    value[2463] = 17'd90901;
    value[2464] = 17'd90894;
    value[2465] = 17'd90887;
    value[2466] = 17'd90879;
    value[2467] = 17'd90872;
    value[2468] = 17'd90865;
    value[2469] = 17'd90858;
    value[2470] = 17'd90850;
    value[2471] = 17'd90843;
    value[2472] = 17'd90836;
    value[2473] = 17'd90828;
    value[2474] = 17'd90821;
    value[2475] = 17'd90814;
    value[2476] = 17'd90807;
    value[2477] = 17'd90799;
    value[2478] = 17'd90792;
    value[2479] = 17'd90785;
    value[2480] = 17'd90777;
    value[2481] = 17'd90770;
    value[2482] = 17'd90763;
    value[2483] = 17'd90755;
    value[2484] = 17'd90748;
    value[2485] = 17'd90741;
    value[2486] = 17'd90733;
    value[2487] = 17'd90726;
    value[2488] = 17'd90719;
    value[2489] = 17'd90711;
    value[2490] = 17'd90704;
    value[2491] = 17'd90697;
    value[2492] = 17'd90689;
    value[2493] = 17'd90682;
    value[2494] = 17'd90674;
    value[2495] = 17'd90667;
    value[2496] = 17'd90660;
    value[2497] = 17'd90652;
    value[2498] = 17'd90645;
    value[2499] = 17'd90638;
    value[2500] = 17'd90630;
    value[2501] = 17'd90623;
    value[2502] = 17'd90616;
    value[2503] = 17'd90608;
    value[2504] = 17'd90601;
    value[2505] = 17'd90593;
    value[2506] = 17'd90586;
    value[2507] = 17'd90579;
    value[2508] = 17'd90571;
    value[2509] = 17'd90564;
    value[2510] = 17'd90556;
    value[2511] = 17'd90549;
    value[2512] = 17'd90542;
    value[2513] = 17'd90534;
    value[2514] = 17'd90527;
    value[2515] = 17'd90519;
    value[2516] = 17'd90512;
    value[2517] = 17'd90504;
    value[2518] = 17'd90497;
    value[2519] = 17'd90490;
    value[2520] = 17'd90482;
    value[2521] = 17'd90475;
    value[2522] = 17'd90467;
    value[2523] = 17'd90460;
    value[2524] = 17'd90452;
    value[2525] = 17'd90445;
    value[2526] = 17'd90438;
    value[2527] = 17'd90430;
    value[2528] = 17'd90423;
    value[2529] = 17'd90415;
    value[2530] = 17'd90408;
    value[2531] = 17'd90400;
    value[2532] = 17'd90393;
    value[2533] = 17'd90385;
    value[2534] = 17'd90378;
    value[2535] = 17'd90370;
    value[2536] = 17'd90363;
    value[2537] = 17'd90355;
    value[2538] = 17'd90348;
    value[2539] = 17'd90341;
    value[2540] = 17'd90333;
    value[2541] = 17'd90326;
    value[2542] = 17'd90318;
    value[2543] = 17'd90311;
    value[2544] = 17'd90303;
    value[2545] = 17'd90296;
    value[2546] = 17'd90288;
    value[2547] = 17'd90281;
    value[2548] = 17'd90273;
    value[2549] = 17'd90266;
    value[2550] = 17'd90258;
    value[2551] = 17'd90251;
    value[2552] = 17'd90243;
    value[2553] = 17'd90235;
    value[2554] = 17'd90228;
    value[2555] = 17'd90220;
    value[2556] = 17'd90213;
    value[2557] = 17'd90205;
    value[2558] = 17'd90198;
    value[2559] = 17'd90190;
    value[2560] = 17'd90183;
    value[2561] = 17'd90175;
    value[2562] = 17'd90168;
    value[2563] = 17'd90160;
    value[2564] = 17'd90153;
    value[2565] = 17'd90145;
    value[2566] = 17'd90137;
    value[2567] = 17'd90130;
    value[2568] = 17'd90122;
    value[2569] = 17'd90115;
    value[2570] = 17'd90107;
    value[2571] = 17'd90100;
    value[2572] = 17'd90092;
    value[2573] = 17'd90084;
    value[2574] = 17'd90077;
    value[2575] = 17'd90069;
    value[2576] = 17'd90062;
    value[2577] = 17'd90054;
    value[2578] = 17'd90047;
    value[2579] = 17'd90039;
    value[2580] = 17'd90031;
    value[2581] = 17'd90024;
    value[2582] = 17'd90016;
    value[2583] = 17'd90009;
    value[2584] = 17'd90001;
    value[2585] = 17'd89993;
    value[2586] = 17'd89986;
    value[2587] = 17'd89978;
    value[2588] = 17'd89971;
    value[2589] = 17'd89963;
    value[2590] = 17'd89955;
    value[2591] = 17'd89948;
    value[2592] = 17'd89940;
    value[2593] = 17'd89932;
    value[2594] = 17'd89925;
    value[2595] = 17'd89917;
    value[2596] = 17'd89909;
    value[2597] = 17'd89902;
    value[2598] = 17'd89894;
    value[2599] = 17'd89887;
    value[2600] = 17'd89879;
    value[2601] = 17'd89871;
    value[2602] = 17'd89864;
    value[2603] = 17'd89856;
    value[2604] = 17'd89848;
    value[2605] = 17'd89841;
    value[2606] = 17'd89833;
    value[2607] = 17'd89825;
    value[2608] = 17'd89818;
    value[2609] = 17'd89810;
    value[2610] = 17'd89802;
    value[2611] = 17'd89795;
    value[2612] = 17'd89787;
    value[2613] = 17'd89779;
    value[2614] = 17'd89772;
    value[2615] = 17'd89764;
    value[2616] = 17'd89756;
    value[2617] = 17'd89748;
    value[2618] = 17'd89741;
    value[2619] = 17'd89733;
    value[2620] = 17'd89725;
    value[2621] = 17'd89718;
    value[2622] = 17'd89710;
    value[2623] = 17'd89702;
    value[2624] = 17'd89694;
    value[2625] = 17'd89687;
    value[2626] = 17'd89679;
    value[2627] = 17'd89671;
    value[2628] = 17'd89664;
    value[2629] = 17'd89656;
    value[2630] = 17'd89648;
    value[2631] = 17'd89640;
    value[2632] = 17'd89633;
    value[2633] = 17'd89625;
    value[2634] = 17'd89617;
    value[2635] = 17'd89609;
    value[2636] = 17'd89602;
    value[2637] = 17'd89594;
    value[2638] = 17'd89586;
    value[2639] = 17'd89578;
    value[2640] = 17'd89571;
    value[2641] = 17'd89563;
    value[2642] = 17'd89555;
    value[2643] = 17'd89547;
    value[2644] = 17'd89540;
    value[2645] = 17'd89532;
    value[2646] = 17'd89524;
    value[2647] = 17'd89516;
    value[2648] = 17'd89509;
    value[2649] = 17'd89501;
    value[2650] = 17'd89493;
    value[2651] = 17'd89485;
    value[2652] = 17'd89477;
    value[2653] = 17'd89470;
    value[2654] = 17'd89462;
    value[2655] = 17'd89454;
    value[2656] = 17'd89446;
    value[2657] = 17'd89438;
    value[2658] = 17'd89431;
    value[2659] = 17'd89423;
    value[2660] = 17'd89415;
    value[2661] = 17'd89407;
    value[2662] = 17'd89399;
    value[2663] = 17'd89391;
    value[2664] = 17'd89384;
    value[2665] = 17'd89376;
    value[2666] = 17'd89368;
    value[2667] = 17'd89360;
    value[2668] = 17'd89352;
    value[2669] = 17'd89344;
    value[2670] = 17'd89337;
    value[2671] = 17'd89329;
    value[2672] = 17'd89321;
    value[2673] = 17'd89313;
    value[2674] = 17'd89305;
    value[2675] = 17'd89297;
    value[2676] = 17'd89290;
    value[2677] = 17'd89282;
    value[2678] = 17'd89274;
    value[2679] = 17'd89266;
    value[2680] = 17'd89258;
    value[2681] = 17'd89250;
    value[2682] = 17'd89242;
    value[2683] = 17'd89234;
    value[2684] = 17'd89227;
    value[2685] = 17'd89219;
    value[2686] = 17'd89211;
    value[2687] = 17'd89203;
    value[2688] = 17'd89195;
    value[2689] = 17'd89187;
    value[2690] = 17'd89179;
    value[2691] = 17'd89171;
    value[2692] = 17'd89163;
    value[2693] = 17'd89156;
    value[2694] = 17'd89148;
    value[2695] = 17'd89140;
    value[2696] = 17'd89132;
    value[2697] = 17'd89124;
    value[2698] = 17'd89116;
    value[2699] = 17'd89108;
    value[2700] = 17'd89100;
    value[2701] = 17'd89092;
    value[2702] = 17'd89084;
    value[2703] = 17'd89076;
    value[2704] = 17'd89068;
    value[2705] = 17'd89061;
    value[2706] = 17'd89053;
    value[2707] = 17'd89045;
    value[2708] = 17'd89037;
    value[2709] = 17'd89029;
    value[2710] = 17'd89021;
    value[2711] = 17'd89013;
    value[2712] = 17'd89005;
    value[2713] = 17'd88997;
    value[2714] = 17'd88989;
    value[2715] = 17'd88981;
    value[2716] = 17'd88973;
    value[2717] = 17'd88965;
    value[2718] = 17'd88957;
    value[2719] = 17'd88949;
    value[2720] = 17'd88941;
    value[2721] = 17'd88933;
    value[2722] = 17'd88925;
    value[2723] = 17'd88917;
    value[2724] = 17'd88909;
    value[2725] = 17'd88901;
    value[2726] = 17'd88893;
    value[2727] = 17'd88885;
    value[2728] = 17'd88877;
    value[2729] = 17'd88869;
    value[2730] = 17'd88861;
    value[2731] = 17'd88853;
    value[2732] = 17'd88845;
    value[2733] = 17'd88837;
    value[2734] = 17'd88829;
    value[2735] = 17'd88821;
    value[2736] = 17'd88813;
    value[2737] = 17'd88805;
    value[2738] = 17'd88797;
    value[2739] = 17'd88789;
    value[2740] = 17'd88781;
    value[2741] = 17'd88773;
    value[2742] = 17'd88765;
    value[2743] = 17'd88757;
    value[2744] = 17'd88749;
    value[2745] = 17'd88741;
    value[2746] = 17'd88733;
    value[2747] = 17'd88725;
    value[2748] = 17'd88717;
    value[2749] = 17'd88709;
    value[2750] = 17'd88701;
    value[2751] = 17'd88693;
    value[2752] = 17'd88684;
    value[2753] = 17'd88676;
    value[2754] = 17'd88668;
    value[2755] = 17'd88660;
    value[2756] = 17'd88652;
    value[2757] = 17'd88644;
    value[2758] = 17'd88636;
    value[2759] = 17'd88628;
    value[2760] = 17'd88620;
    value[2761] = 17'd88612;
    value[2762] = 17'd88604;
    value[2763] = 17'd88596;
    value[2764] = 17'd88587;
    value[2765] = 17'd88579;
    value[2766] = 17'd88571;
    value[2767] = 17'd88563;
    value[2768] = 17'd88555;
    value[2769] = 17'd88547;
    value[2770] = 17'd88539;
    value[2771] = 17'd88531;
    value[2772] = 17'd88523;
    value[2773] = 17'd88515;
    value[2774] = 17'd88506;
    value[2775] = 17'd88498;
    value[2776] = 17'd88490;
    value[2777] = 17'd88482;
    value[2778] = 17'd88474;
    value[2779] = 17'd88466;
    value[2780] = 17'd88458;
    value[2781] = 17'd88449;
    value[2782] = 17'd88441;
    value[2783] = 17'd88433;
    value[2784] = 17'd88425;
    value[2785] = 17'd88417;
    value[2786] = 17'd88409;
    value[2787] = 17'd88401;
    value[2788] = 17'd88392;
    value[2789] = 17'd88384;
    value[2790] = 17'd88376;
    value[2791] = 17'd88368;
    value[2792] = 17'd88360;
    value[2793] = 17'd88352;
    value[2794] = 17'd88343;
    value[2795] = 17'd88335;
    value[2796] = 17'd88327;
    value[2797] = 17'd88319;
    value[2798] = 17'd88311;
    value[2799] = 17'd88302;
    value[2800] = 17'd88294;
    value[2801] = 17'd88286;
    value[2802] = 17'd88278;
    value[2803] = 17'd88270;
    value[2804] = 17'd88261;
    value[2805] = 17'd88253;
    value[2806] = 17'd88245;
    value[2807] = 17'd88237;
    value[2808] = 17'd88229;
    value[2809] = 17'd88220;
    value[2810] = 17'd88212;
    value[2811] = 17'd88204;
    value[2812] = 17'd88196;
    value[2813] = 17'd88188;
    value[2814] = 17'd88179;
    value[2815] = 17'd88171;
    value[2816] = 17'd88163;
    value[2817] = 17'd88155;
    value[2818] = 17'd88146;
    value[2819] = 17'd88138;
    value[2820] = 17'd88130;
    value[2821] = 17'd88122;
    value[2822] = 17'd88113;
    value[2823] = 17'd88105;
    value[2824] = 17'd88097;
    value[2825] = 17'd88089;
    value[2826] = 17'd88080;
    value[2827] = 17'd88072;
    value[2828] = 17'd88064;
    value[2829] = 17'd88056;
    value[2830] = 17'd88047;
    value[2831] = 17'd88039;
    value[2832] = 17'd88031;
    value[2833] = 17'd88022;
    value[2834] = 17'd88014;
    value[2835] = 17'd88006;
    value[2836] = 17'd87998;
    value[2837] = 17'd87989;
    value[2838] = 17'd87981;
    value[2839] = 17'd87973;
    value[2840] = 17'd87964;
    value[2841] = 17'd87956;
    value[2842] = 17'd87948;
    value[2843] = 17'd87939;
    value[2844] = 17'd87931;
    value[2845] = 17'd87923;
    value[2846] = 17'd87915;
    value[2847] = 17'd87906;
    value[2848] = 17'd87898;
    value[2849] = 17'd87890;
    value[2850] = 17'd87881;
    value[2851] = 17'd87873;
    value[2852] = 17'd87865;
    value[2853] = 17'd87856;
    value[2854] = 17'd87848;
    value[2855] = 17'd87840;
    value[2856] = 17'd87831;
    value[2857] = 17'd87823;
    value[2858] = 17'd87815;
    value[2859] = 17'd87806;
    value[2860] = 17'd87798;
    value[2861] = 17'd87789;
    value[2862] = 17'd87781;
    value[2863] = 17'd87773;
    value[2864] = 17'd87764;
    value[2865] = 17'd87756;
    value[2866] = 17'd87748;
    value[2867] = 17'd87739;
    value[2868] = 17'd87731;
    value[2869] = 17'd87723;
    value[2870] = 17'd87714;
    value[2871] = 17'd87706;
    value[2872] = 17'd87697;
    value[2873] = 17'd87689;
    value[2874] = 17'd87681;
    value[2875] = 17'd87672;
    value[2876] = 17'd87664;
    value[2877] = 17'd87655;
    value[2878] = 17'd87647;
    value[2879] = 17'd87639;
    value[2880] = 17'd87630;
    value[2881] = 17'd87622;
    value[2882] = 17'd87613;
    value[2883] = 17'd87605;
    value[2884] = 17'd87597;
    value[2885] = 17'd87588;
    value[2886] = 17'd87580;
    value[2887] = 17'd87571;
    value[2888] = 17'd87563;
    value[2889] = 17'd87554;
    value[2890] = 17'd87546;
    value[2891] = 17'd87538;
    value[2892] = 17'd87529;
    value[2893] = 17'd87521;
    value[2894] = 17'd87512;
    value[2895] = 17'd87504;
    value[2896] = 17'd87495;
    value[2897] = 17'd87487;
    value[2898] = 17'd87478;
    value[2899] = 17'd87470;
    value[2900] = 17'd87461;
    value[2901] = 17'd87453;
    value[2902] = 17'd87445;
    value[2903] = 17'd87436;
    value[2904] = 17'd87428;
    value[2905] = 17'd87419;
    value[2906] = 17'd87411;
    value[2907] = 17'd87402;
    value[2908] = 17'd87394;
    value[2909] = 17'd87385;
    value[2910] = 17'd87377;
    value[2911] = 17'd87368;
    value[2912] = 17'd87360;
    value[2913] = 17'd87351;
    value[2914] = 17'd87343;
    value[2915] = 17'd87334;
    value[2916] = 17'd87326;
    value[2917] = 17'd87317;
    value[2918] = 17'd87309;
    value[2919] = 17'd87300;
    value[2920] = 17'd87292;
    value[2921] = 17'd87283;
    value[2922] = 17'd87275;
    value[2923] = 17'd87266;
    value[2924] = 17'd87258;
    value[2925] = 17'd87249;
    value[2926] = 17'd87241;
    value[2927] = 17'd87232;
    value[2928] = 17'd87224;
    value[2929] = 17'd87215;
    value[2930] = 17'd87206;
    value[2931] = 17'd87198;
    value[2932] = 17'd87189;
    value[2933] = 17'd87181;
    value[2934] = 17'd87172;
    value[2935] = 17'd87164;
    value[2936] = 17'd87155;
    value[2937] = 17'd87147;
    value[2938] = 17'd87138;
    value[2939] = 17'd87129;
    value[2940] = 17'd87121;
    value[2941] = 17'd87112;
    value[2942] = 17'd87104;
    value[2943] = 17'd87095;
    value[2944] = 17'd87087;
    value[2945] = 17'd87078;
    value[2946] = 17'd87069;
    value[2947] = 17'd87061;
    value[2948] = 17'd87052;
    value[2949] = 17'd87044;
    value[2950] = 17'd87035;
    value[2951] = 17'd87026;
    value[2952] = 17'd87018;
    value[2953] = 17'd87009;
    value[2954] = 17'd87001;
    value[2955] = 17'd86992;
    value[2956] = 17'd86983;
    value[2957] = 17'd86975;
    value[2958] = 17'd86966;
    value[2959] = 17'd86958;
    value[2960] = 17'd86949;
    value[2961] = 17'd86940;
    value[2962] = 17'd86932;
    value[2963] = 17'd86923;
    value[2964] = 17'd86914;
    value[2965] = 17'd86906;
    value[2966] = 17'd86897;
    value[2967] = 17'd86889;
    value[2968] = 17'd86880;
    value[2969] = 17'd86871;
    value[2970] = 17'd86863;
    value[2971] = 17'd86854;
    value[2972] = 17'd86845;
    value[2973] = 17'd86837;
    value[2974] = 17'd86828;
    value[2975] = 17'd86819;
    value[2976] = 17'd86811;
    value[2977] = 17'd86802;
    value[2978] = 17'd86793;
    value[2979] = 17'd86785;
    value[2980] = 17'd86776;
    value[2981] = 17'd86767;
    value[2982] = 17'd86759;
    value[2983] = 17'd86750;
    value[2984] = 17'd86741;
    value[2985] = 17'd86733;
    value[2986] = 17'd86724;
    value[2987] = 17'd86715;
    value[2988] = 17'd86707;
    value[2989] = 17'd86698;
    value[2990] = 17'd86689;
    value[2991] = 17'd86680;
    value[2992] = 17'd86672;
    value[2993] = 17'd86663;
    value[2994] = 17'd86654;
    value[2995] = 17'd86646;
    value[2996] = 17'd86637;
    value[2997] = 17'd86628;
    value[2998] = 17'd86619;
    value[2999] = 17'd86611;
    value[3000] = 17'd86602;
    value[3001] = 17'd86593;
    value[3002] = 17'd86585;
    value[3003] = 17'd86576;
    value[3004] = 17'd86567;
    value[3005] = 17'd86558;
    value[3006] = 17'd86550;
    value[3007] = 17'd86541;
    value[3008] = 17'd86532;
    value[3009] = 17'd86523;
    value[3010] = 17'd86515;
    value[3011] = 17'd86506;
    value[3012] = 17'd86497;
    value[3013] = 17'd86488;
    value[3014] = 17'd86480;
    value[3015] = 17'd86471;
    value[3016] = 17'd86462;
    value[3017] = 17'd86453;
    value[3018] = 17'd86445;
    value[3019] = 17'd86436;
    value[3020] = 17'd86427;
    value[3021] = 17'd86418;
    value[3022] = 17'd86409;
    value[3023] = 17'd86401;
    value[3024] = 17'd86392;
    value[3025] = 17'd86383;
    value[3026] = 17'd86374;
    value[3027] = 17'd86365;
    value[3028] = 17'd86357;
    value[3029] = 17'd86348;
    value[3030] = 17'd86339;
    value[3031] = 17'd86330;
    value[3032] = 17'd86321;
    value[3033] = 17'd86313;
    value[3034] = 17'd86304;
    value[3035] = 17'd86295;
    value[3036] = 17'd86286;
    value[3037] = 17'd86277;
    value[3038] = 17'd86269;
    value[3039] = 17'd86260;
    value[3040] = 17'd86251;
    value[3041] = 17'd86242;
    value[3042] = 17'd86233;
    value[3043] = 17'd86224;
    value[3044] = 17'd86216;
    value[3045] = 17'd86207;
    value[3046] = 17'd86198;
    value[3047] = 17'd86189;
    value[3048] = 17'd86180;
    value[3049] = 17'd86171;
    value[3050] = 17'd86162;
    value[3051] = 17'd86154;
    value[3052] = 17'd86145;
    value[3053] = 17'd86136;
    value[3054] = 17'd86127;
    value[3055] = 17'd86118;
    value[3056] = 17'd86109;
    value[3057] = 17'd86100;
    value[3058] = 17'd86091;
    value[3059] = 17'd86083;
    value[3060] = 17'd86074;
    value[3061] = 17'd86065;
    value[3062] = 17'd86056;
    value[3063] = 17'd86047;
    value[3064] = 17'd86038;
    value[3065] = 17'd86029;
    value[3066] = 17'd86020;
    value[3067] = 17'd86011;
    value[3068] = 17'd86003;
    value[3069] = 17'd85994;
    value[3070] = 17'd85985;
    value[3071] = 17'd85976;
    value[3072] = 17'd85967;
    value[3073] = 17'd85958;
    value[3074] = 17'd85949;
    value[3075] = 17'd85940;
    value[3076] = 17'd85931;
    value[3077] = 17'd85922;
    value[3078] = 17'd85913;
    value[3079] = 17'd85904;
    value[3080] = 17'd85895;
    value[3081] = 17'd85887;
    value[3082] = 17'd85878;
    value[3083] = 17'd85869;
    value[3084] = 17'd85860;
    value[3085] = 17'd85851;
    value[3086] = 17'd85842;
    value[3087] = 17'd85833;
    value[3088] = 17'd85824;
    value[3089] = 17'd85815;
    value[3090] = 17'd85806;
    value[3091] = 17'd85797;
    value[3092] = 17'd85788;
    value[3093] = 17'd85779;
    value[3094] = 17'd85770;
    value[3095] = 17'd85761;
    value[3096] = 17'd85752;
    value[3097] = 17'd85743;
    value[3098] = 17'd85734;
    value[3099] = 17'd85725;
    value[3100] = 17'd85716;
    value[3101] = 17'd85707;
    value[3102] = 17'd85698;
    value[3103] = 17'd85689;
    value[3104] = 17'd85680;
    value[3105] = 17'd85671;
    value[3106] = 17'd85662;
    value[3107] = 17'd85653;
    value[3108] = 17'd85644;
    value[3109] = 17'd85635;
    value[3110] = 17'd85626;
    value[3111] = 17'd85617;
    value[3112] = 17'd85608;
    value[3113] = 17'd85599;
    value[3114] = 17'd85590;
    value[3115] = 17'd85581;
    value[3116] = 17'd85572;
    value[3117] = 17'd85563;
    value[3118] = 17'd85554;
    value[3119] = 17'd85545;
    value[3120] = 17'd85536;
    value[3121] = 17'd85527;
    value[3122] = 17'd85518;
    value[3123] = 17'd85509;
    value[3124] = 17'd85500;
    value[3125] = 17'd85491;
    value[3126] = 17'd85482;
    value[3127] = 17'd85473;
    value[3128] = 17'd85464;
    value[3129] = 17'd85454;
    value[3130] = 17'd85445;
    value[3131] = 17'd85436;
    value[3132] = 17'd85427;
    value[3133] = 17'd85418;
    value[3134] = 17'd85409;
    value[3135] = 17'd85400;
    value[3136] = 17'd85391;
    value[3137] = 17'd85382;
    value[3138] = 17'd85373;
    value[3139] = 17'd85364;
    value[3140] = 17'd85355;
    value[3141] = 17'd85345;
    value[3142] = 17'd85336;
    value[3143] = 17'd85327;
    value[3144] = 17'd85318;
    value[3145] = 17'd85309;
    value[3146] = 17'd85300;
    value[3147] = 17'd85291;
    value[3148] = 17'd85282;
    value[3149] = 17'd85273;
    value[3150] = 17'd85264;
    value[3151] = 17'd85254;
    value[3152] = 17'd85245;
    value[3153] = 17'd85236;
    value[3154] = 17'd85227;
    value[3155] = 17'd85218;
    value[3156] = 17'd85209;
    value[3157] = 17'd85200;
    value[3158] = 17'd85190;
    value[3159] = 17'd85181;
    value[3160] = 17'd85172;
    value[3161] = 17'd85163;
    value[3162] = 17'd85154;
    value[3163] = 17'd85145;
    value[3164] = 17'd85136;
    value[3165] = 17'd85126;
    value[3166] = 17'd85117;
    value[3167] = 17'd85108;
    value[3168] = 17'd85099;
    value[3169] = 17'd85090;
    value[3170] = 17'd85081;
    value[3171] = 17'd85071;
    value[3172] = 17'd85062;
    value[3173] = 17'd85053;
    value[3174] = 17'd85044;
    value[3175] = 17'd85035;
    value[3176] = 17'd85026;
    value[3177] = 17'd85016;
    value[3178] = 17'd85007;
    value[3179] = 17'd84998;
    value[3180] = 17'd84989;
    value[3181] = 17'd84980;
    value[3182] = 17'd84970;
    value[3183] = 17'd84961;
    value[3184] = 17'd84952;
    value[3185] = 17'd84943;
    value[3186] = 17'd84934;
    value[3187] = 17'd84924;
    value[3188] = 17'd84915;
    value[3189] = 17'd84906;
    value[3190] = 17'd84897;
    value[3191] = 17'd84887;
    value[3192] = 17'd84878;
    value[3193] = 17'd84869;
    value[3194] = 17'd84860;
    value[3195] = 17'd84851;
    value[3196] = 17'd84841;
    value[3197] = 17'd84832;
    value[3198] = 17'd84823;
    value[3199] = 17'd84814;
    value[3200] = 17'd84804;
    value[3201] = 17'd84795;
    value[3202] = 17'd84786;
    value[3203] = 17'd84777;
    value[3204] = 17'd84767;
    value[3205] = 17'd84758;
    value[3206] = 17'd84749;
    value[3207] = 17'd84740;
    value[3208] = 17'd84730;
    value[3209] = 17'd84721;
    value[3210] = 17'd84712;
    value[3211] = 17'd84702;
    value[3212] = 17'd84693;
    value[3213] = 17'd84684;
    value[3214] = 17'd84675;
    value[3215] = 17'd84665;
    value[3216] = 17'd84656;
    value[3217] = 17'd84647;
    value[3218] = 17'd84637;
    value[3219] = 17'd84628;
    value[3220] = 17'd84619;
    value[3221] = 17'd84610;
    value[3222] = 17'd84600;
    value[3223] = 17'd84591;
    value[3224] = 17'd84582;
    value[3225] = 17'd84572;
    value[3226] = 17'd84563;
    value[3227] = 17'd84554;
    value[3228] = 17'd84544;
    value[3229] = 17'd84535;
    value[3230] = 17'd84526;
    value[3231] = 17'd84516;
    value[3232] = 17'd84507;
    value[3233] = 17'd84498;
    value[3234] = 17'd84488;
    value[3235] = 17'd84479;
    value[3236] = 17'd84470;
    value[3237] = 17'd84460;
    value[3238] = 17'd84451;
    value[3239] = 17'd84442;
    value[3240] = 17'd84432;
    value[3241] = 17'd84423;
    value[3242] = 17'd84414;
    value[3243] = 17'd84404;
    value[3244] = 17'd84395;
    value[3245] = 17'd84386;
    value[3246] = 17'd84376;
    value[3247] = 17'd84367;
    value[3248] = 17'd84357;
    value[3249] = 17'd84348;
    value[3250] = 17'd84339;
    value[3251] = 17'd84329;
    value[3252] = 17'd84320;
    value[3253] = 17'd84311;
    value[3254] = 17'd84301;
    value[3255] = 17'd84292;
    value[3256] = 17'd84282;
    value[3257] = 17'd84273;
    value[3258] = 17'd84264;
    value[3259] = 17'd84254;
    value[3260] = 17'd84245;
    value[3261] = 17'd84235;
    value[3262] = 17'd84226;
    value[3263] = 17'd84217;
    value[3264] = 17'd84207;
    value[3265] = 17'd84198;
    value[3266] = 17'd84188;
    value[3267] = 17'd84179;
    value[3268] = 17'd84169;
    value[3269] = 17'd84160;
    value[3270] = 17'd84151;
    value[3271] = 17'd84141;
    value[3272] = 17'd84132;
    value[3273] = 17'd84122;
    value[3274] = 17'd84113;
    value[3275] = 17'd84103;
    value[3276] = 17'd84094;
    value[3277] = 17'd84085;
    value[3278] = 17'd84075;
    value[3279] = 17'd84066;
    value[3280] = 17'd84056;
    value[3281] = 17'd84047;
    value[3282] = 17'd84037;
    value[3283] = 17'd84028;
    value[3284] = 17'd84018;
    value[3285] = 17'd84009;
    value[3286] = 17'd83999;
    value[3287] = 17'd83990;
    value[3288] = 17'd83980;
    value[3289] = 17'd83971;
    value[3290] = 17'd83961;
    value[3291] = 17'd83952;
    value[3292] = 17'd83943;
    value[3293] = 17'd83933;
    value[3294] = 17'd83924;
    value[3295] = 17'd83914;
    value[3296] = 17'd83905;
    value[3297] = 17'd83895;
    value[3298] = 17'd83886;
    value[3299] = 17'd83876;
    value[3300] = 17'd83867;
    value[3301] = 17'd83857;
    value[3302] = 17'd83848;
    value[3303] = 17'd83838;
    value[3304] = 17'd83829;
    value[3305] = 17'd83819;
    value[3306] = 17'd83809;
    value[3307] = 17'd83800;
    value[3308] = 17'd83790;
    value[3309] = 17'd83781;
    value[3310] = 17'd83771;
    value[3311] = 17'd83762;
    value[3312] = 17'd83752;
    value[3313] = 17'd83743;
    value[3314] = 17'd83733;
    value[3315] = 17'd83724;
    value[3316] = 17'd83714;
    value[3317] = 17'd83705;
    value[3318] = 17'd83695;
    value[3319] = 17'd83685;
    value[3320] = 17'd83676;
    value[3321] = 17'd83666;
    value[3322] = 17'd83657;
    value[3323] = 17'd83647;
    value[3324] = 17'd83638;
    value[3325] = 17'd83628;
    value[3326] = 17'd83619;
    value[3327] = 17'd83609;
    value[3328] = 17'd83599;
    value[3329] = 17'd83590;
    value[3330] = 17'd83580;
    value[3331] = 17'd83571;
    value[3332] = 17'd83561;
    value[3333] = 17'd83551;
    value[3334] = 17'd83542;
    value[3335] = 17'd83532;
    value[3336] = 17'd83523;
    value[3337] = 17'd83513;
    value[3338] = 17'd83504;
    value[3339] = 17'd83494;
    value[3340] = 17'd83484;
    value[3341] = 17'd83475;
    value[3342] = 17'd83465;
    value[3343] = 17'd83455;
    value[3344] = 17'd83446;
    value[3345] = 17'd83436;
    value[3346] = 17'd83427;
    value[3347] = 17'd83417;
    value[3348] = 17'd83407;
    value[3349] = 17'd83398;
    value[3350] = 17'd83388;
    value[3351] = 17'd83378;
    value[3352] = 17'd83369;
    value[3353] = 17'd83359;
    value[3354] = 17'd83350;
    value[3355] = 17'd83340;
    value[3356] = 17'd83330;
    value[3357] = 17'd83321;
    value[3358] = 17'd83311;
    value[3359] = 17'd83301;
    value[3360] = 17'd83292;
    value[3361] = 17'd83282;
    value[3362] = 17'd83272;
    value[3363] = 17'd83263;
    value[3364] = 17'd83253;
    value[3365] = 17'd83243;
    value[3366] = 17'd83234;
    value[3367] = 17'd83224;
    value[3368] = 17'd83214;
    value[3369] = 17'd83205;
    value[3370] = 17'd83195;
    value[3371] = 17'd83185;
    value[3372] = 17'd83176;
    value[3373] = 17'd83166;
    value[3374] = 17'd83156;
    value[3375] = 17'd83146;
    value[3376] = 17'd83137;
    value[3377] = 17'd83127;
    value[3378] = 17'd83117;
    value[3379] = 17'd83108;
    value[3380] = 17'd83098;
    value[3381] = 17'd83088;
    value[3382] = 17'd83079;
    value[3383] = 17'd83069;
    value[3384] = 17'd83059;
    value[3385] = 17'd83049;
    value[3386] = 17'd83040;
    value[3387] = 17'd83030;
    value[3388] = 17'd83020;
    value[3389] = 17'd83010;
    value[3390] = 17'd83001;
    value[3391] = 17'd82991;
    value[3392] = 17'd82981;
    value[3393] = 17'd82972;
    value[3394] = 17'd82962;
    value[3395] = 17'd82952;
    value[3396] = 17'd82942;
    value[3397] = 17'd82933;
    value[3398] = 17'd82923;
    value[3399] = 17'd82913;
    value[3400] = 17'd82903;
    value[3401] = 17'd82894;
    value[3402] = 17'd82884;
    value[3403] = 17'd82874;
    value[3404] = 17'd82864;
    value[3405] = 17'd82854;
    value[3406] = 17'd82845;
    value[3407] = 17'd82835;
    value[3408] = 17'd82825;
    value[3409] = 17'd82815;
    value[3410] = 17'd82806;
    value[3411] = 17'd82796;
    value[3412] = 17'd82786;
    value[3413] = 17'd82776;
    value[3414] = 17'd82766;
    value[3415] = 17'd82757;
    value[3416] = 17'd82747;
    value[3417] = 17'd82737;
    value[3418] = 17'd82727;
    value[3419] = 17'd82717;
    value[3420] = 17'd82708;
    value[3421] = 17'd82698;
    value[3422] = 17'd82688;
    value[3423] = 17'd82678;
    value[3424] = 17'd82668;
    value[3425] = 17'd82658;
    value[3426] = 17'd82649;
    value[3427] = 17'd82639;
    value[3428] = 17'd82629;
    value[3429] = 17'd82619;
    value[3430] = 17'd82609;
    value[3431] = 17'd82599;
    value[3432] = 17'd82590;
    value[3433] = 17'd82580;
    value[3434] = 17'd82570;
    value[3435] = 17'd82560;
    value[3436] = 17'd82550;
    value[3437] = 17'd82540;
    value[3438] = 17'd82531;
    value[3439] = 17'd82521;
    value[3440] = 17'd82511;
    value[3441] = 17'd82501;
    value[3442] = 17'd82491;
    value[3443] = 17'd82481;
    value[3444] = 17'd82471;
    value[3445] = 17'd82462;
    value[3446] = 17'd82452;
    value[3447] = 17'd82442;
    value[3448] = 17'd82432;
    value[3449] = 17'd82422;
    value[3450] = 17'd82412;
    value[3451] = 17'd82402;
    value[3452] = 17'd82392;
    value[3453] = 17'd82382;
    value[3454] = 17'd82373;
    value[3455] = 17'd82363;
    value[3456] = 17'd82353;
    value[3457] = 17'd82343;
    value[3458] = 17'd82333;
    value[3459] = 17'd82323;
    value[3460] = 17'd82313;
    value[3461] = 17'd82303;
    value[3462] = 17'd82293;
    value[3463] = 17'd82283;
    value[3464] = 17'd82273;
    value[3465] = 17'd82264;
    value[3466] = 17'd82254;
    value[3467] = 17'd82244;
    value[3468] = 17'd82234;
    value[3469] = 17'd82224;
    value[3470] = 17'd82214;
    value[3471] = 17'd82204;
    value[3472] = 17'd82194;
    value[3473] = 17'd82184;
    value[3474] = 17'd82174;
    value[3475] = 17'd82164;
    value[3476] = 17'd82154;
    value[3477] = 17'd82144;
    value[3478] = 17'd82134;
    value[3479] = 17'd82124;
    value[3480] = 17'd82114;
    value[3481] = 17'd82104;
    value[3482] = 17'd82094;
    value[3483] = 17'd82085;
    value[3484] = 17'd82075;
    value[3485] = 17'd82065;
    value[3486] = 17'd82055;
    value[3487] = 17'd82045;
    value[3488] = 17'd82035;
    value[3489] = 17'd82025;
    value[3490] = 17'd82015;
    value[3491] = 17'd82005;
    value[3492] = 17'd81995;
    value[3493] = 17'd81985;
    value[3494] = 17'd81975;
    value[3495] = 17'd81965;
    value[3496] = 17'd81955;
    value[3497] = 17'd81945;
    value[3498] = 17'd81935;
    value[3499] = 17'd81925;
    value[3500] = 17'd81915;
    value[3501] = 17'd81905;
    value[3502] = 17'd81895;
    value[3503] = 17'd81885;
    value[3504] = 17'd81875;
    value[3505] = 17'd81865;
    value[3506] = 17'd81855;
    value[3507] = 17'd81845;
    value[3508] = 17'd81835;
    value[3509] = 17'd81825;
    value[3510] = 17'd81814;
    value[3511] = 17'd81804;
    value[3512] = 17'd81794;
    value[3513] = 17'd81784;
    value[3514] = 17'd81774;
    value[3515] = 17'd81764;
    value[3516] = 17'd81754;
    value[3517] = 17'd81744;
    value[3518] = 17'd81734;
    value[3519] = 17'd81724;
    value[3520] = 17'd81714;
    value[3521] = 17'd81704;
    value[3522] = 17'd81694;
    value[3523] = 17'd81684;
    value[3524] = 17'd81674;
    value[3525] = 17'd81664;
    value[3526] = 17'd81654;
    value[3527] = 17'd81644;
    value[3528] = 17'd81633;
    value[3529] = 17'd81623;
    value[3530] = 17'd81613;
    value[3531] = 17'd81603;
    value[3532] = 17'd81593;
    value[3533] = 17'd81583;
    value[3534] = 17'd81573;
    value[3535] = 17'd81563;
    value[3536] = 17'd81553;
    value[3537] = 17'd81543;
    value[3538] = 17'd81532;
    value[3539] = 17'd81522;
    value[3540] = 17'd81512;
    value[3541] = 17'd81502;
    value[3542] = 17'd81492;
    value[3543] = 17'd81482;
    value[3544] = 17'd81472;
    value[3545] = 17'd81462;
    value[3546] = 17'd81452;
    value[3547] = 17'd81441;
    value[3548] = 17'd81431;
    value[3549] = 17'd81421;
    value[3550] = 17'd81411;
    value[3551] = 17'd81401;
    value[3552] = 17'd81391;
    value[3553] = 17'd81381;
    value[3554] = 17'd81370;
    value[3555] = 17'd81360;
    value[3556] = 17'd81350;
    value[3557] = 17'd81340;
    value[3558] = 17'd81330;
    value[3559] = 17'd81320;
    value[3560] = 17'd81310;
    value[3561] = 17'd81299;
    value[3562] = 17'd81289;
    value[3563] = 17'd81279;
    value[3564] = 17'd81269;
    value[3565] = 17'd81259;
    value[3566] = 17'd81249;
    value[3567] = 17'd81238;
    value[3568] = 17'd81228;
    value[3569] = 17'd81218;
    value[3570] = 17'd81208;
    value[3571] = 17'd81198;
    value[3572] = 17'd81187;
    value[3573] = 17'd81177;
    value[3574] = 17'd81167;
    value[3575] = 17'd81157;
    value[3576] = 17'd81147;
    value[3577] = 17'd81137;
    value[3578] = 17'd81126;
    value[3579] = 17'd81116;
    value[3580] = 17'd81106;
    value[3581] = 17'd81096;
    value[3582] = 17'd81085;
    value[3583] = 17'd81075;
    value[3584] = 17'd81065;
    value[3585] = 17'd81055;
    value[3586] = 17'd81045;
    value[3587] = 17'd81034;
    value[3588] = 17'd81024;
    value[3589] = 17'd81014;
    value[3590] = 17'd81004;
    value[3591] = 17'd80993;
    value[3592] = 17'd80983;
    value[3593] = 17'd80973;
    value[3594] = 17'd80963;
    value[3595] = 17'd80952;
    value[3596] = 17'd80942;
    value[3597] = 17'd80932;
    value[3598] = 17'd80922;
    value[3599] = 17'd80911;
    value[3600] = 17'd80901;
    value[3601] = 17'd80891;
    value[3602] = 17'd80881;
    value[3603] = 17'd80870;
    value[3604] = 17'd80860;
    value[3605] = 17'd80850;
    value[3606] = 17'd80840;
    value[3607] = 17'd80829;
    value[3608] = 17'd80819;
    value[3609] = 17'd80809;
    value[3610] = 17'd80798;
    value[3611] = 17'd80788;
    value[3612] = 17'd80778;
    value[3613] = 17'd80768;
    value[3614] = 17'd80757;
    value[3615] = 17'd80747;
    value[3616] = 17'd80737;
    value[3617] = 17'd80726;
    value[3618] = 17'd80716;
    value[3619] = 17'd80706;
    value[3620] = 17'd80696;
    value[3621] = 17'd80685;
    value[3622] = 17'd80675;
    value[3623] = 17'd80665;
    value[3624] = 17'd80654;
    value[3625] = 17'd80644;
    value[3626] = 17'd80634;
    value[3627] = 17'd80623;
    value[3628] = 17'd80613;
    value[3629] = 17'd80603;
    value[3630] = 17'd80592;
    value[3631] = 17'd80582;
    value[3632] = 17'd80572;
    value[3633] = 17'd80561;
    value[3634] = 17'd80551;
    value[3635] = 17'd80541;
    value[3636] = 17'd80530;
    value[3637] = 17'd80520;
    value[3638] = 17'd80510;
    value[3639] = 17'd80499;
    value[3640] = 17'd80489;
    value[3641] = 17'd80479;
    value[3642] = 17'd80468;
    value[3643] = 17'd80458;
    value[3644] = 17'd80447;
    value[3645] = 17'd80437;
    value[3646] = 17'd80427;
    value[3647] = 17'd80416;
    value[3648] = 17'd80406;
    value[3649] = 17'd80396;
    value[3650] = 17'd80385;
    value[3651] = 17'd80375;
    value[3652] = 17'd80364;
    value[3653] = 17'd80354;
    value[3654] = 17'd80344;
    value[3655] = 17'd80333;
    value[3656] = 17'd80323;
    value[3657] = 17'd80312;
    value[3658] = 17'd80302;
    value[3659] = 17'd80292;
    value[3660] = 17'd80281;
    value[3661] = 17'd80271;
    value[3662] = 17'd80260;
    value[3663] = 17'd80250;
    value[3664] = 17'd80240;
    value[3665] = 17'd80229;
    value[3666] = 17'd80219;
    value[3667] = 17'd80208;
    value[3668] = 17'd80198;
    value[3669] = 17'd80187;
    value[3670] = 17'd80177;
    value[3671] = 17'd80167;
    value[3672] = 17'd80156;
    value[3673] = 17'd80146;
    value[3674] = 17'd80135;
    value[3675] = 17'd80125;
    value[3676] = 17'd80114;
    value[3677] = 17'd80104;
    value[3678] = 17'd80094;
    value[3679] = 17'd80083;
    value[3680] = 17'd80073;
    value[3681] = 17'd80062;
    value[3682] = 17'd80052;
    value[3683] = 17'd80041;
    value[3684] = 17'd80031;
    value[3685] = 17'd80020;
    value[3686] = 17'd80010;
    value[3687] = 17'd79999;
    value[3688] = 17'd79989;
    value[3689] = 17'd79978;
    value[3690] = 17'd79968;
    value[3691] = 17'd79957;
    value[3692] = 17'd79947;
    value[3693] = 17'd79937;
    value[3694] = 17'd79926;
    value[3695] = 17'd79916;
    value[3696] = 17'd79905;
    value[3697] = 17'd79895;
    value[3698] = 17'd79884;
    value[3699] = 17'd79874;
    value[3700] = 17'd79863;
    value[3701] = 17'd79853;
    value[3702] = 17'd79842;
    value[3703] = 17'd79832;
    value[3704] = 17'd79821;
    value[3705] = 17'd79811;
    value[3706] = 17'd79800;
    value[3707] = 17'd79789;
    value[3708] = 17'd79779;
    value[3709] = 17'd79768;
    value[3710] = 17'd79758;
    value[3711] = 17'd79747;
    value[3712] = 17'd79737;
    value[3713] = 17'd79726;
    value[3714] = 17'd79716;
    value[3715] = 17'd79705;
    value[3716] = 17'd79695;
    value[3717] = 17'd79684;
    value[3718] = 17'd79674;
    value[3719] = 17'd79663;
    value[3720] = 17'd79652;
    value[3721] = 17'd79642;
    value[3722] = 17'd79631;
    value[3723] = 17'd79621;
    value[3724] = 17'd79610;
    value[3725] = 17'd79600;
    value[3726] = 17'd79589;
    value[3727] = 17'd79579;
    value[3728] = 17'd79568;
    value[3729] = 17'd79557;
    value[3730] = 17'd79547;
    value[3731] = 17'd79536;
    value[3732] = 17'd79526;
    value[3733] = 17'd79515;
    value[3734] = 17'd79505;
    value[3735] = 17'd79494;
    value[3736] = 17'd79483;
    value[3737] = 17'd79473;
    value[3738] = 17'd79462;
    value[3739] = 17'd79452;
    value[3740] = 17'd79441;
    value[3741] = 17'd79430;
    value[3742] = 17'd79420;
    value[3743] = 17'd79409;
    value[3744] = 17'd79399;
    value[3745] = 17'd79388;
    value[3746] = 17'd79377;
    value[3747] = 17'd79367;
    value[3748] = 17'd79356;
    value[3749] = 17'd79345;
    value[3750] = 17'd79335;
    value[3751] = 17'd79324;
    value[3752] = 17'd79314;
    value[3753] = 17'd79303;
    value[3754] = 17'd79292;
    value[3755] = 17'd79282;
    value[3756] = 17'd79271;
    value[3757] = 17'd79260;
    value[3758] = 17'd79250;
    value[3759] = 17'd79239;
    value[3760] = 17'd79228;
    value[3761] = 17'd79218;
    value[3762] = 17'd79207;
    value[3763] = 17'd79197;
    value[3764] = 17'd79186;
    value[3765] = 17'd79175;
    value[3766] = 17'd79165;
    value[3767] = 17'd79154;
    value[3768] = 17'd79143;
    value[3769] = 17'd79133;
    value[3770] = 17'd79122;
    value[3771] = 17'd79111;
    value[3772] = 17'd79101;
    value[3773] = 17'd79090;
    value[3774] = 17'd79079;
    value[3775] = 17'd79068;
    value[3776] = 17'd79058;
    value[3777] = 17'd79047;
    value[3778] = 17'd79036;
    value[3779] = 17'd79026;
    value[3780] = 17'd79015;
    value[3781] = 17'd79004;
    value[3782] = 17'd78994;
    value[3783] = 17'd78983;
    value[3784] = 17'd78972;
    value[3785] = 17'd78961;
    value[3786] = 17'd78951;
    value[3787] = 17'd78940;
    value[3788] = 17'd78929;
    value[3789] = 17'd78919;
    value[3790] = 17'd78908;
    value[3791] = 17'd78897;
    value[3792] = 17'd78886;
    value[3793] = 17'd78876;
    value[3794] = 17'd78865;
    value[3795] = 17'd78854;
    value[3796] = 17'd78844;
    value[3797] = 17'd78833;
    value[3798] = 17'd78822;
    value[3799] = 17'd78811;
    value[3800] = 17'd78801;
    value[3801] = 17'd78790;
    value[3802] = 17'd78779;
    value[3803] = 17'd78768;
    value[3804] = 17'd78758;
    value[3805] = 17'd78747;
    value[3806] = 17'd78736;
    value[3807] = 17'd78725;
    value[3808] = 17'd78715;
    value[3809] = 17'd78704;
    value[3810] = 17'd78693;
    value[3811] = 17'd78682;
    value[3812] = 17'd78671;
    value[3813] = 17'd78661;
    value[3814] = 17'd78650;
    value[3815] = 17'd78639;
    value[3816] = 17'd78628;
    value[3817] = 17'd78618;
    value[3818] = 17'd78607;
    value[3819] = 17'd78596;
    value[3820] = 17'd78585;
    value[3821] = 17'd78574;
    value[3822] = 17'd78564;
    value[3823] = 17'd78553;
    value[3824] = 17'd78542;
    value[3825] = 17'd78531;
    value[3826] = 17'd78520;
    value[3827] = 17'd78510;
    value[3828] = 17'd78499;
    value[3829] = 17'd78488;
    value[3830] = 17'd78477;
    value[3831] = 17'd78466;
    value[3832] = 17'd78456;
    value[3833] = 17'd78445;
    value[3834] = 17'd78434;
    value[3835] = 17'd78423;
    value[3836] = 17'd78412;
    value[3837] = 17'd78401;
    value[3838] = 17'd78391;
    value[3839] = 17'd78380;
    value[3840] = 17'd78369;
    value[3841] = 17'd78358;
    value[3842] = 17'd78347;
    value[3843] = 17'd78336;
    value[3844] = 17'd78325;
    value[3845] = 17'd78315;
    value[3846] = 17'd78304;
    value[3847] = 17'd78293;
    value[3848] = 17'd78282;
    value[3849] = 17'd78271;
    value[3850] = 17'd78260;
    value[3851] = 17'd78249;
    value[3852] = 17'd78239;
    value[3853] = 17'd78228;
    value[3854] = 17'd78217;
    value[3855] = 17'd78206;
    value[3856] = 17'd78195;
    value[3857] = 17'd78184;
    value[3858] = 17'd78173;
    value[3859] = 17'd78162;
    value[3860] = 17'd78152;
    value[3861] = 17'd78141;
    value[3862] = 17'd78130;
    value[3863] = 17'd78119;
    value[3864] = 17'd78108;
    value[3865] = 17'd78097;
    value[3866] = 17'd78086;
    value[3867] = 17'd78075;
    value[3868] = 17'd78064;
    value[3869] = 17'd78053;
    value[3870] = 17'd78043;
    value[3871] = 17'd78032;
    value[3872] = 17'd78021;
    value[3873] = 17'd78010;
    value[3874] = 17'd77999;
    value[3875] = 17'd77988;
    value[3876] = 17'd77977;
    value[3877] = 17'd77966;
    value[3878] = 17'd77955;
    value[3879] = 17'd77944;
    value[3880] = 17'd77933;
    value[3881] = 17'd77922;
    value[3882] = 17'd77911;
    value[3883] = 17'd77900;
    value[3884] = 17'd77890;
    value[3885] = 17'd77879;
    value[3886] = 17'd77868;
    value[3887] = 17'd77857;
    value[3888] = 17'd77846;
    value[3889] = 17'd77835;
    value[3890] = 17'd77824;
    value[3891] = 17'd77813;
    value[3892] = 17'd77802;
    value[3893] = 17'd77791;
    value[3894] = 17'd77780;
    value[3895] = 17'd77769;
    value[3896] = 17'd77758;
    value[3897] = 17'd77747;
    value[3898] = 17'd77736;
    value[3899] = 17'd77725;
    value[3900] = 17'd77714;
    value[3901] = 17'd77703;
    value[3902] = 17'd77692;
    value[3903] = 17'd77681;
    value[3904] = 17'd77670;
    value[3905] = 17'd77659;
    value[3906] = 17'd77648;
    value[3907] = 17'd77637;
    value[3908] = 17'd77626;
    value[3909] = 17'd77615;
    value[3910] = 17'd77604;
    value[3911] = 17'd77593;
    value[3912] = 17'd77582;
    value[3913] = 17'd77571;
    value[3914] = 17'd77560;
    value[3915] = 17'd77549;
    value[3916] = 17'd77538;
    value[3917] = 17'd77527;
    value[3918] = 17'd77516;
    value[3919] = 17'd77505;
    value[3920] = 17'd77494;
    value[3921] = 17'd77483;
    value[3922] = 17'd77472;
    value[3923] = 17'd77461;
    value[3924] = 17'd77450;
    value[3925] = 17'd77439;
    value[3926] = 17'd77428;
    value[3927] = 17'd77417;
    value[3928] = 17'd77406;
    value[3929] = 17'd77395;
    value[3930] = 17'd77384;
    value[3931] = 17'd77372;
    value[3932] = 17'd77361;
    value[3933] = 17'd77350;
    value[3934] = 17'd77339;
    value[3935] = 17'd77328;
    value[3936] = 17'd77317;
    value[3937] = 17'd77306;
    value[3938] = 17'd77295;
    value[3939] = 17'd77284;
    value[3940] = 17'd77273;
    value[3941] = 17'd77262;
    value[3942] = 17'd77251;
    value[3943] = 17'd77240;
    value[3944] = 17'd77229;
    value[3945] = 17'd77217;
    value[3946] = 17'd77206;
    value[3947] = 17'd77195;
    value[3948] = 17'd77184;
    value[3949] = 17'd77173;
    value[3950] = 17'd77162;
    value[3951] = 17'd77151;
    value[3952] = 17'd77140;
    value[3953] = 17'd77129;
    value[3954] = 17'd77118;
    value[3955] = 17'd77106;
    value[3956] = 17'd77095;
    value[3957] = 17'd77084;
    value[3958] = 17'd77073;
    value[3959] = 17'd77062;
    value[3960] = 17'd77051;
    value[3961] = 17'd77040;
    value[3962] = 17'd77029;
    value[3963] = 17'd77017;
    value[3964] = 17'd77006;
    value[3965] = 17'd76995;
    value[3966] = 17'd76984;
    value[3967] = 17'd76973;
    value[3968] = 17'd76962;
    value[3969] = 17'd76951;
    value[3970] = 17'd76939;
    value[3971] = 17'd76928;
    value[3972] = 17'd76917;
    value[3973] = 17'd76906;
    value[3974] = 17'd76895;
    value[3975] = 17'd76884;
    value[3976] = 17'd76873;
    value[3977] = 17'd76861;
    value[3978] = 17'd76850;
    value[3979] = 17'd76839;
    value[3980] = 17'd76828;
    value[3981] = 17'd76817;
    value[3982] = 17'd76806;
    value[3983] = 17'd76794;
    value[3984] = 17'd76783;
    value[3985] = 17'd76772;
    value[3986] = 17'd76761;
    value[3987] = 17'd76750;
    value[3988] = 17'd76738;
    value[3989] = 17'd76727;
    value[3990] = 17'd76716;
    value[3991] = 17'd76705;
    value[3992] = 17'd76694;
    value[3993] = 17'd76682;
    value[3994] = 17'd76671;
    value[3995] = 17'd76660;
    value[3996] = 17'd76649;
    value[3997] = 17'd76638;
    value[3998] = 17'd76626;
    value[3999] = 17'd76615;
    value[4000] = 17'd76604;
    value[4001] = 17'd76593;
    value[4002] = 17'd76582;
    value[4003] = 17'd76570;
    value[4004] = 17'd76559;
    value[4005] = 17'd76548;
    value[4006] = 17'd76537;
    value[4007] = 17'd76525;
    value[4008] = 17'd76514;
    value[4009] = 17'd76503;
    value[4010] = 17'd76492;
    value[4011] = 17'd76480;
    value[4012] = 17'd76469;
    value[4013] = 17'd76458;
    value[4014] = 17'd76447;
    value[4015] = 17'd76435;
    value[4016] = 17'd76424;
    value[4017] = 17'd76413;
    value[4018] = 17'd76402;
    value[4019] = 17'd76390;
    value[4020] = 17'd76379;
    value[4021] = 17'd76368;
    value[4022] = 17'd76357;
    value[4023] = 17'd76345;
    value[4024] = 17'd76334;
    value[4025] = 17'd76323;
    value[4026] = 17'd76311;
    value[4027] = 17'd76300;
    value[4028] = 17'd76289;
    value[4029] = 17'd76278;
    value[4030] = 17'd76266;
    value[4031] = 17'd76255;
    value[4032] = 17'd76244;
    value[4033] = 17'd76232;
    value[4034] = 17'd76221;
    value[4035] = 17'd76210;
    value[4036] = 17'd76199;
    value[4037] = 17'd76187;
    value[4038] = 17'd76176;
    value[4039] = 17'd76165;
    value[4040] = 17'd76153;
    value[4041] = 17'd76142;
    value[4042] = 17'd76131;
    value[4043] = 17'd76119;
    value[4044] = 17'd76108;
    value[4045] = 17'd76097;
    value[4046] = 17'd76085;
    value[4047] = 17'd76074;
    value[4048] = 17'd76063;
    value[4049] = 17'd76051;
    value[4050] = 17'd76040;
    value[4051] = 17'd76029;
    value[4052] = 17'd76017;
    value[4053] = 17'd76006;
    value[4054] = 17'd75995;
    value[4055] = 17'd75983;
    value[4056] = 17'd75972;
    value[4057] = 17'd75961;
    value[4058] = 17'd75949;
    value[4059] = 17'd75938;
    value[4060] = 17'd75927;
    value[4061] = 17'd75915;
    value[4062] = 17'd75904;
    value[4063] = 17'd75893;
    value[4064] = 17'd75881;
    value[4065] = 17'd75870;
    value[4066] = 17'd75858;
    value[4067] = 17'd75847;
    value[4068] = 17'd75836;
    value[4069] = 17'd75824;
    value[4070] = 17'd75813;
    value[4071] = 17'd75802;
    value[4072] = 17'd75790;
    value[4073] = 17'd75779;
    value[4074] = 17'd75767;
    value[4075] = 17'd75756;
    value[4076] = 17'd75745;
    value[4077] = 17'd75733;
    value[4078] = 17'd75722;
    value[4079] = 17'd75710;
    value[4080] = 17'd75699;
    value[4081] = 17'd75688;
    value[4082] = 17'd75676;
    value[4083] = 17'd75665;
    value[4084] = 17'd75653;
    value[4085] = 17'd75642;
    value[4086] = 17'd75631;
    value[4087] = 17'd75619;
    value[4088] = 17'd75608;
    value[4089] = 17'd75596;
    value[4090] = 17'd75585;
    value[4091] = 17'd75573;
    value[4092] = 17'd75562;
    value[4093] = 17'd75551;
    value[4094] = 17'd75539;
    value[4095] = 17'd75528;
    value[4096] = 17'd75516;
    value[4097] = 17'd75505;
    value[4098] = 17'd75493;
    value[4099] = 17'd75482;
    value[4100] = 17'd75470;
    value[4101] = 17'd75459;
    value[4102] = 17'd75448;
    value[4103] = 17'd75436;
    value[4104] = 17'd75425;
    value[4105] = 17'd75413;
    value[4106] = 17'd75402;
    value[4107] = 17'd75390;
    value[4108] = 17'd75379;
    value[4109] = 17'd75367;
    value[4110] = 17'd75356;
    value[4111] = 17'd75344;
    value[4112] = 17'd75333;
    value[4113] = 17'd75321;
    value[4114] = 17'd75310;
    value[4115] = 17'd75298;
    value[4116] = 17'd75287;
    value[4117] = 17'd75275;
    value[4118] = 17'd75264;
    value[4119] = 17'd75252;
    value[4120] = 17'd75241;
    value[4121] = 17'd75229;
    value[4122] = 17'd75218;
    value[4123] = 17'd75206;
    value[4124] = 17'd75195;
    value[4125] = 17'd75183;
    value[4126] = 17'd75172;
    value[4127] = 17'd75160;
    value[4128] = 17'd75149;
    value[4129] = 17'd75137;
    value[4130] = 17'd75126;
    value[4131] = 17'd75114;
    value[4132] = 17'd75103;
    value[4133] = 17'd75091;
    value[4134] = 17'd75080;
    value[4135] = 17'd75068;
    value[4136] = 17'd75057;
    value[4137] = 17'd75045;
    value[4138] = 17'd75034;
    value[4139] = 17'd75022;
    value[4140] = 17'd75011;
    value[4141] = 17'd74999;
    value[4142] = 17'd74988;
    value[4143] = 17'd74976;
    value[4144] = 17'd74964;
    value[4145] = 17'd74953;
    value[4146] = 17'd74941;
    value[4147] = 17'd74930;
    value[4148] = 17'd74918;
    value[4149] = 17'd74907;
    value[4150] = 17'd74895;
    value[4151] = 17'd74884;
    value[4152] = 17'd74872;
    value[4153] = 17'd74860;
    value[4154] = 17'd74849;
    value[4155] = 17'd74837;
    value[4156] = 17'd74826;
    value[4157] = 17'd74814;
    value[4158] = 17'd74802;
    value[4159] = 17'd74791;
    value[4160] = 17'd74779;
    value[4161] = 17'd74768;
    value[4162] = 17'd74756;
    value[4163] = 17'd74745;
    value[4164] = 17'd74733;
    value[4165] = 17'd74721;
    value[4166] = 17'd74710;
    value[4167] = 17'd74698;
    value[4168] = 17'd74687;
    value[4169] = 17'd74675;
    value[4170] = 17'd74663;
    value[4171] = 17'd74652;
    value[4172] = 17'd74640;
    value[4173] = 17'd74628;
    value[4174] = 17'd74617;
    value[4175] = 17'd74605;
    value[4176] = 17'd74594;
    value[4177] = 17'd74582;
    value[4178] = 17'd74570;
    value[4179] = 17'd74559;
    value[4180] = 17'd74547;
    value[4181] = 17'd74535;
    value[4182] = 17'd74524;
    value[4183] = 17'd74512;
    value[4184] = 17'd74501;
    value[4185] = 17'd74489;
    value[4186] = 17'd74477;
    value[4187] = 17'd74466;
    value[4188] = 17'd74454;
    value[4189] = 17'd74442;
    value[4190] = 17'd74431;
    value[4191] = 17'd74419;
    value[4192] = 17'd74407;
    value[4193] = 17'd74396;
    value[4194] = 17'd74384;
    value[4195] = 17'd74372;
    value[4196] = 17'd74361;
    value[4197] = 17'd74349;
    value[4198] = 17'd74337;
    value[4199] = 17'd74326;
    value[4200] = 17'd74314;
    value[4201] = 17'd74302;
    value[4202] = 17'd74291;
    value[4203] = 17'd74279;
    value[4204] = 17'd74267;
    value[4205] = 17'd74256;
    value[4206] = 17'd74244;
    value[4207] = 17'd74232;
    value[4208] = 17'd74220;
    value[4209] = 17'd74209;
    value[4210] = 17'd74197;
    value[4211] = 17'd74185;
    value[4212] = 17'd74174;
    value[4213] = 17'd74162;
    value[4214] = 17'd74150;
    value[4215] = 17'd74139;
    value[4216] = 17'd74127;
    value[4217] = 17'd74115;
    value[4218] = 17'd74103;
    value[4219] = 17'd74092;
    value[4220] = 17'd74080;
    value[4221] = 17'd74068;
    value[4222] = 17'd74057;
    value[4223] = 17'd74045;
    value[4224] = 17'd74033;
    value[4225] = 17'd74021;
    value[4226] = 17'd74010;
    value[4227] = 17'd73998;
    value[4228] = 17'd73986;
    value[4229] = 17'd73974;
    value[4230] = 17'd73963;
    value[4231] = 17'd73951;
    value[4232] = 17'd73939;
    value[4233] = 17'd73927;
    value[4234] = 17'd73916;
    value[4235] = 17'd73904;
    value[4236] = 17'd73892;
    value[4237] = 17'd73880;
    value[4238] = 17'd73869;
    value[4239] = 17'd73857;
    value[4240] = 17'd73845;
    value[4241] = 17'd73833;
    value[4242] = 17'd73821;
    value[4243] = 17'd73810;
    value[4244] = 17'd73798;
    value[4245] = 17'd73786;
    value[4246] = 17'd73774;
    value[4247] = 17'd73763;
    value[4248] = 17'd73751;
    value[4249] = 17'd73739;
    value[4250] = 17'd73727;
    value[4251] = 17'd73715;
    value[4252] = 17'd73704;
    value[4253] = 17'd73692;
    value[4254] = 17'd73680;
    value[4255] = 17'd73668;
    value[4256] = 17'd73656;
    value[4257] = 17'd73645;
    value[4258] = 17'd73633;
    value[4259] = 17'd73621;
    value[4260] = 17'd73609;
    value[4261] = 17'd73597;
    value[4262] = 17'd73586;
    value[4263] = 17'd73574;
    value[4264] = 17'd73562;
    value[4265] = 17'd73550;
    value[4266] = 17'd73538;
    value[4267] = 17'd73526;
    value[4268] = 17'd73515;
    value[4269] = 17'd73503;
    value[4270] = 17'd73491;
    value[4271] = 17'd73479;
    value[4272] = 17'd73467;
    value[4273] = 17'd73455;
    value[4274] = 17'd73444;
    value[4275] = 17'd73432;
    value[4276] = 17'd73420;
    value[4277] = 17'd73408;
    value[4278] = 17'd73396;
    value[4279] = 17'd73384;
    value[4280] = 17'd73372;
    value[4281] = 17'd73361;
    value[4282] = 17'd73349;
    value[4283] = 17'd73337;
    value[4284] = 17'd73325;
    value[4285] = 17'd73313;
    value[4286] = 17'd73301;
    value[4287] = 17'd73289;
    value[4288] = 17'd73278;
    value[4289] = 17'd73266;
    value[4290] = 17'd73254;
    value[4291] = 17'd73242;
    value[4292] = 17'd73230;
    value[4293] = 17'd73218;
    value[4294] = 17'd73206;
    value[4295] = 17'd73194;
    value[4296] = 17'd73182;
    value[4297] = 17'd73171;
    value[4298] = 17'd73159;
    value[4299] = 17'd73147;
    value[4300] = 17'd73135;
    value[4301] = 17'd73123;
    value[4302] = 17'd73111;
    value[4303] = 17'd73099;
    value[4304] = 17'd73087;
    value[4305] = 17'd73075;
    value[4306] = 17'd73063;
    value[4307] = 17'd73051;
    value[4308] = 17'd73040;
    value[4309] = 17'd73028;
    value[4310] = 17'd73016;
    value[4311] = 17'd73004;
    value[4312] = 17'd72992;
    value[4313] = 17'd72980;
    value[4314] = 17'd72968;
    value[4315] = 17'd72956;
    value[4316] = 17'd72944;
    value[4317] = 17'd72932;
    value[4318] = 17'd72920;
    value[4319] = 17'd72908;
    value[4320] = 17'd72896;
    value[4321] = 17'd72884;
    value[4322] = 17'd72872;
    value[4323] = 17'd72861;
    value[4324] = 17'd72849;
    value[4325] = 17'd72837;
    value[4326] = 17'd72825;
    value[4327] = 17'd72813;
    value[4328] = 17'd72801;
    value[4329] = 17'd72789;
    value[4330] = 17'd72777;
    value[4331] = 17'd72765;
    value[4332] = 17'd72753;
    value[4333] = 17'd72741;
    value[4334] = 17'd72729;
    value[4335] = 17'd72717;
    value[4336] = 17'd72705;
    value[4337] = 17'd72693;
    value[4338] = 17'd72681;
    value[4339] = 17'd72669;
    value[4340] = 17'd72657;
    value[4341] = 17'd72645;
    value[4342] = 17'd72633;
    value[4343] = 17'd72621;
    value[4344] = 17'd72609;
    value[4345] = 17'd72597;
    value[4346] = 17'd72585;
    value[4347] = 17'd72573;
    value[4348] = 17'd72561;
    value[4349] = 17'd72549;
    value[4350] = 17'd72537;
    value[4351] = 17'd72525;
    value[4352] = 17'd72513;
    value[4353] = 17'd72501;
    value[4354] = 17'd72489;
    value[4355] = 17'd72477;
    value[4356] = 17'd72465;
    value[4357] = 17'd72453;
    value[4358] = 17'd72441;
    value[4359] = 17'd72429;
    value[4360] = 17'd72417;
    value[4361] = 17'd72405;
    value[4362] = 17'd72393;
    value[4363] = 17'd72381;
    value[4364] = 17'd72369;
    value[4365] = 17'd72356;
    value[4366] = 17'd72344;
    value[4367] = 17'd72332;
    value[4368] = 17'd72320;
    value[4369] = 17'd72308;
    value[4370] = 17'd72296;
    value[4371] = 17'd72284;
    value[4372] = 17'd72272;
    value[4373] = 17'd72260;
    value[4374] = 17'd72248;
    value[4375] = 17'd72236;
    value[4376] = 17'd72224;
    value[4377] = 17'd72212;
    value[4378] = 17'd72200;
    value[4379] = 17'd72188;
    value[4380] = 17'd72176;
    value[4381] = 17'd72163;
    value[4382] = 17'd72151;
    value[4383] = 17'd72139;
    value[4384] = 17'd72127;
    value[4385] = 17'd72115;
    value[4386] = 17'd72103;
    value[4387] = 17'd72091;
    value[4388] = 17'd72079;
    value[4389] = 17'd72067;
    value[4390] = 17'd72055;
    value[4391] = 17'd72043;
    value[4392] = 17'd72030;
    value[4393] = 17'd72018;
    value[4394] = 17'd72006;
    value[4395] = 17'd71994;
    value[4396] = 17'd71982;
    value[4397] = 17'd71970;
    value[4398] = 17'd71958;
    value[4399] = 17'd71946;
    value[4400] = 17'd71933;
    value[4401] = 17'd71921;
    value[4402] = 17'd71909;
    value[4403] = 17'd71897;
    value[4404] = 17'd71885;
    value[4405] = 17'd71873;
    value[4406] = 17'd71861;
    value[4407] = 17'd71849;
    value[4408] = 17'd71836;
    value[4409] = 17'd71824;
    value[4410] = 17'd71812;
    value[4411] = 17'd71800;
    value[4412] = 17'd71788;
    value[4413] = 17'd71776;
    value[4414] = 17'd71764;
    value[4415] = 17'd71751;
    value[4416] = 17'd71739;
    value[4417] = 17'd71727;
    value[4418] = 17'd71715;
    value[4419] = 17'd71703;
    value[4420] = 17'd71691;
    value[4421] = 17'd71678;
    value[4422] = 17'd71666;
    value[4423] = 17'd71654;
    value[4424] = 17'd71642;
    value[4425] = 17'd71630;
    value[4426] = 17'd71618;
    value[4427] = 17'd71605;
    value[4428] = 17'd71593;
    value[4429] = 17'd71581;
    value[4430] = 17'd71569;
    value[4431] = 17'd71557;
    value[4432] = 17'd71544;
    value[4433] = 17'd71532;
    value[4434] = 17'd71520;
    value[4435] = 17'd71508;
    value[4436] = 17'd71496;
    value[4437] = 17'd71483;
    value[4438] = 17'd71471;
    value[4439] = 17'd71459;
    value[4440] = 17'd71447;
    value[4441] = 17'd71435;
    value[4442] = 17'd71422;
    value[4443] = 17'd71410;
    value[4444] = 17'd71398;
    value[4445] = 17'd71386;
    value[4446] = 17'd71373;
    value[4447] = 17'd71361;
    value[4448] = 17'd71349;
    value[4449] = 17'd71337;
    value[4450] = 17'd71325;
    value[4451] = 17'd71312;
    value[4452] = 17'd71300;
    value[4453] = 17'd71288;
    value[4454] = 17'd71276;
    value[4455] = 17'd71263;
    value[4456] = 17'd71251;
    value[4457] = 17'd71239;
    value[4458] = 17'd71227;
    value[4459] = 17'd71214;
    value[4460] = 17'd71202;
    value[4461] = 17'd71190;
    value[4462] = 17'd71178;
    value[4463] = 17'd71165;
    value[4464] = 17'd71153;
    value[4465] = 17'd71141;
    value[4466] = 17'd71129;
    value[4467] = 17'd71116;
    value[4468] = 17'd71104;
    value[4469] = 17'd71092;
    value[4470] = 17'd71079;
    value[4471] = 17'd71067;
    value[4472] = 17'd71055;
    value[4473] = 17'd71043;
    value[4474] = 17'd71030;
    value[4475] = 17'd71018;
    value[4476] = 17'd71006;
    value[4477] = 17'd70993;
    value[4478] = 17'd70981;
    value[4479] = 17'd70969;
    value[4480] = 17'd70957;
    value[4481] = 17'd70944;
    value[4482] = 17'd70932;
    value[4483] = 17'd70920;
    value[4484] = 17'd70907;
    value[4485] = 17'd70895;
    value[4486] = 17'd70883;
    value[4487] = 17'd70870;
    value[4488] = 17'd70858;
    value[4489] = 17'd70846;
    value[4490] = 17'd70833;
    value[4491] = 17'd70821;
    value[4492] = 17'd70809;
    value[4493] = 17'd70797;
    value[4494] = 17'd70784;
    value[4495] = 17'd70772;
    value[4496] = 17'd70760;
    value[4497] = 17'd70747;
    value[4498] = 17'd70735;
    value[4499] = 17'd70723;
    value[4500] = 17'd70710;
    value[4501] = 17'd70698;
    value[4502] = 17'd70685;
    value[4503] = 17'd70673;
    value[4504] = 17'd70661;
    value[4505] = 17'd70648;
    value[4506] = 17'd70636;
    value[4507] = 17'd70624;
    value[4508] = 17'd70611;
    value[4509] = 17'd70599;
    value[4510] = 17'd70587;
    value[4511] = 17'd70574;
    value[4512] = 17'd70562;
    value[4513] = 17'd70550;
    value[4514] = 17'd70537;
    value[4515] = 17'd70525;
    value[4516] = 17'd70512;
    value[4517] = 17'd70500;
    value[4518] = 17'd70488;
    value[4519] = 17'd70475;
    value[4520] = 17'd70463;
    value[4521] = 17'd70451;
    value[4522] = 17'd70438;
    value[4523] = 17'd70426;
    value[4524] = 17'd70413;
    value[4525] = 17'd70401;
    value[4526] = 17'd70389;
    value[4527] = 17'd70376;
    value[4528] = 17'd70364;
    value[4529] = 17'd70351;
    value[4530] = 17'd70339;
    value[4531] = 17'd70327;
    value[4532] = 17'd70314;
    value[4533] = 17'd70302;
    value[4534] = 17'd70289;
    value[4535] = 17'd70277;
    value[4536] = 17'd70265;
    value[4537] = 17'd70252;
    value[4538] = 17'd70240;
    value[4539] = 17'd70227;
    value[4540] = 17'd70215;
    value[4541] = 17'd70202;
    value[4542] = 17'd70190;
    value[4543] = 17'd70178;
    value[4544] = 17'd70165;
    value[4545] = 17'd70153;
    value[4546] = 17'd70140;
    value[4547] = 17'd70128;
    value[4548] = 17'd70115;
    value[4549] = 17'd70103;
    value[4550] = 17'd70090;
    value[4551] = 17'd70078;
    value[4552] = 17'd70066;
    value[4553] = 17'd70053;
    value[4554] = 17'd70041;
    value[4555] = 17'd70028;
    value[4556] = 17'd70016;
    value[4557] = 17'd70003;
    value[4558] = 17'd69991;
    value[4559] = 17'd69978;
    value[4560] = 17'd69966;
    value[4561] = 17'd69953;
    value[4562] = 17'd69941;
    value[4563] = 17'd69928;
    value[4564] = 17'd69916;
    value[4565] = 17'd69903;
    value[4566] = 17'd69891;
    value[4567] = 17'd69878;
    value[4568] = 17'd69866;
    value[4569] = 17'd69854;
    value[4570] = 17'd69841;
    value[4571] = 17'd69829;
    value[4572] = 17'd69816;
    value[4573] = 17'd69804;
    value[4574] = 17'd69791;
    value[4575] = 17'd69779;
    value[4576] = 17'd69766;
    value[4577] = 17'd69754;
    value[4578] = 17'd69741;
    value[4579] = 17'd69729;
    value[4580] = 17'd69716;
    value[4581] = 17'd69704;
    value[4582] = 17'd69691;
    value[4583] = 17'd69678;
    value[4584] = 17'd69666;
    value[4585] = 17'd69653;
    value[4586] = 17'd69641;
    value[4587] = 17'd69628;
    value[4588] = 17'd69616;
    value[4589] = 17'd69603;
    value[4590] = 17'd69591;
    value[4591] = 17'd69578;
    value[4592] = 17'd69566;
    value[4593] = 17'd69553;
    value[4594] = 17'd69541;
    value[4595] = 17'd69528;
    value[4596] = 17'd69516;
    value[4597] = 17'd69503;
    value[4598] = 17'd69490;
    value[4599] = 17'd69478;
    value[4600] = 17'd69465;
    value[4601] = 17'd69453;
    value[4602] = 17'd69440;
    value[4603] = 17'd69428;
    value[4604] = 17'd69415;
    value[4605] = 17'd69403;
    value[4606] = 17'd69390;
    value[4607] = 17'd69377;
    value[4608] = 17'd69365;
    value[4609] = 17'd69352;
    value[4610] = 17'd69340;
    value[4611] = 17'd69327;
    value[4612] = 17'd69315;
    value[4613] = 17'd69302;
    value[4614] = 17'd69289;
    value[4615] = 17'd69277;
    value[4616] = 17'd69264;
    value[4617] = 17'd69252;
    value[4618] = 17'd69239;
    value[4619] = 17'd69226;
    value[4620] = 17'd69214;
    value[4621] = 17'd69201;
    value[4622] = 17'd69189;
    value[4623] = 17'd69176;
    value[4624] = 17'd69163;
    value[4625] = 17'd69151;
    value[4626] = 17'd69138;
    value[4627] = 17'd69126;
    value[4628] = 17'd69113;
    value[4629] = 17'd69100;
    value[4630] = 17'd69088;
    value[4631] = 17'd69075;
    value[4632] = 17'd69063;
    value[4633] = 17'd69050;
    value[4634] = 17'd69037;
    value[4635] = 17'd69025;
    value[4636] = 17'd69012;
    value[4637] = 17'd68999;
    value[4638] = 17'd68987;
    value[4639] = 17'd68974;
    value[4640] = 17'd68961;
    value[4641] = 17'd68949;
    value[4642] = 17'd68936;
    value[4643] = 17'd68924;
    value[4644] = 17'd68911;
    value[4645] = 17'd68898;
    value[4646] = 17'd68886;
    value[4647] = 17'd68873;
    value[4648] = 17'd68860;
    value[4649] = 17'd68848;
    value[4650] = 17'd68835;
    value[4651] = 17'd68822;
    value[4652] = 17'd68810;
    value[4653] = 17'd68797;
    value[4654] = 17'd68784;
    value[4655] = 17'd68772;
    value[4656] = 17'd68759;
    value[4657] = 17'd68746;
    value[4658] = 17'd68734;
    value[4659] = 17'd68721;
    value[4660] = 17'd68708;
    value[4661] = 17'd68696;
    value[4662] = 17'd68683;
    value[4663] = 17'd68670;
    value[4664] = 17'd68658;
    value[4665] = 17'd68645;
    value[4666] = 17'd68632;
    value[4667] = 17'd68619;
    value[4668] = 17'd68607;
    value[4669] = 17'd68594;
    value[4670] = 17'd68581;
    value[4671] = 17'd68569;
    value[4672] = 17'd68556;
    value[4673] = 17'd68543;
    value[4674] = 17'd68531;
    value[4675] = 17'd68518;
    value[4676] = 17'd68505;
    value[4677] = 17'd68492;
    value[4678] = 17'd68480;
    value[4679] = 17'd68467;
    value[4680] = 17'd68454;
    value[4681] = 17'd68441;
    value[4682] = 17'd68429;
    value[4683] = 17'd68416;
    value[4684] = 17'd68403;
    value[4685] = 17'd68391;
    value[4686] = 17'd68378;
    value[4687] = 17'd68365;
    value[4688] = 17'd68352;
    value[4689] = 17'd68340;
    value[4690] = 17'd68327;
    value[4691] = 17'd68314;
    value[4692] = 17'd68301;
    value[4693] = 17'd68289;
    value[4694] = 17'd68276;
    value[4695] = 17'd68263;
    value[4696] = 17'd68250;
    value[4697] = 17'd68238;
    value[4698] = 17'd68225;
    value[4699] = 17'd68212;
    value[4700] = 17'd68199;
    value[4701] = 17'd68187;
    value[4702] = 17'd68174;
    value[4703] = 17'd68161;
    value[4704] = 17'd68148;
    value[4705] = 17'd68135;
    value[4706] = 17'd68123;
    value[4707] = 17'd68110;
    value[4708] = 17'd68097;
    value[4709] = 17'd68084;
    value[4710] = 17'd68072;
    value[4711] = 17'd68059;
    value[4712] = 17'd68046;
    value[4713] = 17'd68033;
    value[4714] = 17'd68020;
    value[4715] = 17'd68008;
    value[4716] = 17'd67995;
    value[4717] = 17'd67982;
    value[4718] = 17'd67969;
    value[4719] = 17'd67956;
    value[4720] = 17'd67944;
    value[4721] = 17'd67931;
    value[4722] = 17'd67918;
    value[4723] = 17'd67905;
    value[4724] = 17'd67892;
    value[4725] = 17'd67880;
    value[4726] = 17'd67867;
    value[4727] = 17'd67854;
    value[4728] = 17'd67841;
    value[4729] = 17'd67828;
    value[4730] = 17'd67815;
    value[4731] = 17'd67803;
    value[4732] = 17'd67790;
    value[4733] = 17'd67777;
    value[4734] = 17'd67764;
    value[4735] = 17'd67751;
    value[4736] = 17'd67738;
    value[4737] = 17'd67726;
    value[4738] = 17'd67713;
    value[4739] = 17'd67700;
    value[4740] = 17'd67687;
    value[4741] = 17'd67674;
    value[4742] = 17'd67661;
    value[4743] = 17'd67649;
    value[4744] = 17'd67636;
    value[4745] = 17'd67623;
    value[4746] = 17'd67610;
    value[4747] = 17'd67597;
    value[4748] = 17'd67584;
    value[4749] = 17'd67571;
    value[4750] = 17'd67559;
    value[4751] = 17'd67546;
    value[4752] = 17'd67533;
    value[4753] = 17'd67520;
    value[4754] = 17'd67507;
    value[4755] = 17'd67494;
    value[4756] = 17'd67481;
    value[4757] = 17'd67468;
    value[4758] = 17'd67456;
    value[4759] = 17'd67443;
    value[4760] = 17'd67430;
    value[4761] = 17'd67417;
    value[4762] = 17'd67404;
    value[4763] = 17'd67391;
    value[4764] = 17'd67378;
    value[4765] = 17'd67365;
    value[4766] = 17'd67352;
    value[4767] = 17'd67339;
    value[4768] = 17'd67327;
    value[4769] = 17'd67314;
    value[4770] = 17'd67301;
    value[4771] = 17'd67288;
    value[4772] = 17'd67275;
    value[4773] = 17'd67262;
    value[4774] = 17'd67249;
    value[4775] = 17'd67236;
    value[4776] = 17'd67223;
    value[4777] = 17'd67210;
    value[4778] = 17'd67197;
    value[4779] = 17'd67184;
    value[4780] = 17'd67172;
    value[4781] = 17'd67159;
    value[4782] = 17'd67146;
    value[4783] = 17'd67133;
    value[4784] = 17'd67120;
    value[4785] = 17'd67107;
    value[4786] = 17'd67094;
    value[4787] = 17'd67081;
    value[4788] = 17'd67068;
    value[4789] = 17'd67055;
    value[4790] = 17'd67042;
    value[4791] = 17'd67029;
    value[4792] = 17'd67016;
    value[4793] = 17'd67003;
    value[4794] = 17'd66990;
    value[4795] = 17'd66977;
    value[4796] = 17'd66964;
    value[4797] = 17'd66951;
    value[4798] = 17'd66939;
    value[4799] = 17'd66926;
    value[4800] = 17'd66913;
    value[4801] = 17'd66900;
    value[4802] = 17'd66887;
    value[4803] = 17'd66874;
    value[4804] = 17'd66861;
    value[4805] = 17'd66848;
    value[4806] = 17'd66835;
    value[4807] = 17'd66822;
    value[4808] = 17'd66809;
    value[4809] = 17'd66796;
    value[4810] = 17'd66783;
    value[4811] = 17'd66770;
    value[4812] = 17'd66757;
    value[4813] = 17'd66744;
    value[4814] = 17'd66731;
    value[4815] = 17'd66718;
    value[4816] = 17'd66705;
    value[4817] = 17'd66692;
    value[4818] = 17'd66679;
    value[4819] = 17'd66666;
    value[4820] = 17'd66653;
    value[4821] = 17'd66640;
    value[4822] = 17'd66627;
    value[4823] = 17'd66614;
    value[4824] = 17'd66601;
    value[4825] = 17'd66588;
    value[4826] = 17'd66575;
    value[4827] = 17'd66562;
    value[4828] = 17'd66549;
    value[4829] = 17'd66536;
    value[4830] = 17'd66523;
    value[4831] = 17'd66510;
    value[4832] = 17'd66496;
    value[4833] = 17'd66483;
    value[4834] = 17'd66470;
    value[4835] = 17'd66457;
    value[4836] = 17'd66444;
    value[4837] = 17'd66431;
    value[4838] = 17'd66418;
    value[4839] = 17'd66405;
    value[4840] = 17'd66392;
    value[4841] = 17'd66379;
    value[4842] = 17'd66366;
    value[4843] = 17'd66353;
    value[4844] = 17'd66340;
    value[4845] = 17'd66327;
    value[4846] = 17'd66314;
    value[4847] = 17'd66301;
    value[4848] = 17'd66288;
    value[4849] = 17'd66275;
    value[4850] = 17'd66262;
    value[4851] = 17'd66248;
    value[4852] = 17'd66235;
    value[4853] = 17'd66222;
    value[4854] = 17'd66209;
    value[4855] = 17'd66196;
    value[4856] = 17'd66183;
    value[4857] = 17'd66170;
    value[4858] = 17'd66157;
    value[4859] = 17'd66144;
    value[4860] = 17'd66131;
    value[4861] = 17'd66118;
    value[4862] = 17'd66105;
    value[4863] = 17'd66091;
    value[4864] = 17'd66078;
    value[4865] = 17'd66065;
    value[4866] = 17'd66052;
    value[4867] = 17'd66039;
    value[4868] = 17'd66026;
    value[4869] = 17'd66013;
    value[4870] = 17'd66000;
    value[4871] = 17'd65987;
    value[4872] = 17'd65973;
    value[4873] = 17'd65960;
    value[4874] = 17'd65947;
    value[4875] = 17'd65934;
    value[4876] = 17'd65921;
    value[4877] = 17'd65908;
    value[4878] = 17'd65895;
    value[4879] = 17'd65882;
    value[4880] = 17'd65868;
    value[4881] = 17'd65855;
    value[4882] = 17'd65842;
    value[4883] = 17'd65829;
    value[4884] = 17'd65816;
    value[4885] = 17'd65803;
    value[4886] = 17'd65790;
    value[4887] = 17'd65776;
    value[4888] = 17'd65763;
    value[4889] = 17'd65750;
    value[4890] = 17'd65737;
    value[4891] = 17'd65724;
    value[4892] = 17'd65711;
    value[4893] = 17'd65698;
    value[4894] = 17'd65684;
    value[4895] = 17'd65671;
    value[4896] = 17'd65658;
    value[4897] = 17'd65645;
    value[4898] = 17'd65632;
    value[4899] = 17'd65619;
    value[4900] = 17'd65605;
    value[4901] = 17'd65592;
    value[4902] = 17'd65579;
    value[4903] = 17'd65566;
    value[4904] = 17'd65553;
    value[4905] = 17'd65540;
    value[4906] = 17'd65526;
    value[4907] = 17'd65513;
    value[4908] = 17'd65500;
    value[4909] = 17'd65487;
    value[4910] = 17'd65474;
    value[4911] = 17'd65460;
    value[4912] = 17'd65447;
    value[4913] = 17'd65434;
    value[4914] = 17'd65421;
    value[4915] = 17'd65408;
    value[4916] = 17'd65394;
    value[4917] = 17'd65381;
    value[4918] = 17'd65368;
    value[4919] = 17'd65355;
    value[4920] = 17'd65342;
    value[4921] = 17'd65328;
    value[4922] = 17'd65315;
    value[4923] = 17'd65302;
    value[4924] = 17'd65289;
    value[4925] = 17'd65275;
    value[4926] = 17'd65262;
    value[4927] = 17'd65249;
    value[4928] = 17'd65236;
    value[4929] = 17'd65223;
    value[4930] = 17'd65209;
    value[4931] = 17'd65196;
    value[4932] = 17'd65183;
    value[4933] = 17'd65170;
    value[4934] = 17'd65156;
    value[4935] = 17'd65143;
    value[4936] = 17'd65130;
    value[4937] = 17'd65117;
    value[4938] = 17'd65103;
    value[4939] = 17'd65090;
    value[4940] = 17'd65077;
    value[4941] = 17'd65064;
    value[4942] = 17'd65050;
    value[4943] = 17'd65037;
    value[4944] = 17'd65024;
    value[4945] = 17'd65011;
    value[4946] = 17'd64997;
    value[4947] = 17'd64984;
    value[4948] = 17'd64971;
    value[4949] = 17'd64958;
    value[4950] = 17'd64944;
    value[4951] = 17'd64931;
    value[4952] = 17'd64918;
    value[4953] = 17'd64904;
    value[4954] = 17'd64891;
    value[4955] = 17'd64878;
    value[4956] = 17'd64865;
    value[4957] = 17'd64851;
    value[4958] = 17'd64838;
    value[4959] = 17'd64825;
    value[4960] = 17'd64811;
    value[4961] = 17'd64798;
    value[4962] = 17'd64785;
    value[4963] = 17'd64772;
    value[4964] = 17'd64758;
    value[4965] = 17'd64745;
    value[4966] = 17'd64732;
    value[4967] = 17'd64718;
    value[4968] = 17'd64705;
    value[4969] = 17'd64692;
    value[4970] = 17'd64678;
    value[4971] = 17'd64665;
    value[4972] = 17'd64652;
    value[4973] = 17'd64639;
    value[4974] = 17'd64625;
    value[4975] = 17'd64612;
    value[4976] = 17'd64599;
    value[4977] = 17'd64585;
    value[4978] = 17'd64572;
    value[4979] = 17'd64559;
    value[4980] = 17'd64545;
    value[4981] = 17'd64532;
    value[4982] = 17'd64519;
    value[4983] = 17'd64505;
    value[4984] = 17'd64492;
    value[4985] = 17'd64479;
    value[4986] = 17'd64465;
    value[4987] = 17'd64452;
    value[4988] = 17'd64439;
    value[4989] = 17'd64425;
    value[4990] = 17'd64412;
    value[4991] = 17'd64399;
    value[4992] = 17'd64385;
    value[4993] = 17'd64372;
    value[4994] = 17'd64358;
    value[4995] = 17'd64345;
    value[4996] = 17'd64332;
    value[4997] = 17'd64318;
    value[4998] = 17'd64305;
    value[4999] = 17'd64292;
    value[5000] = 17'd64278;
    value[5001] = 17'd64265;
    value[5002] = 17'd64252;
    value[5003] = 17'd64238;
    value[5004] = 17'd64225;
    value[5005] = 17'd64211;
    value[5006] = 17'd64198;
    value[5007] = 17'd64185;
    value[5008] = 17'd64171;
    value[5009] = 17'd64158;
    value[5010] = 17'd64144;
    value[5011] = 17'd64131;
    value[5012] = 17'd64118;
    value[5013] = 17'd64104;
    value[5014] = 17'd64091;
    value[5015] = 17'd64077;
    value[5016] = 17'd64064;
    value[5017] = 17'd64051;
    value[5018] = 17'd64037;
    value[5019] = 17'd64024;
    value[5020] = 17'd64010;
    value[5021] = 17'd63997;
    value[5022] = 17'd63984;
    value[5023] = 17'd63970;
    value[5024] = 17'd63957;
    value[5025] = 17'd63943;
    value[5026] = 17'd63930;
    value[5027] = 17'd63917;
    value[5028] = 17'd63903;
    value[5029] = 17'd63890;
    value[5030] = 17'd63876;
    value[5031] = 17'd63863;
    value[5032] = 17'd63849;
    value[5033] = 17'd63836;
    value[5034] = 17'd63823;
    value[5035] = 17'd63809;
    value[5036] = 17'd63796;
    value[5037] = 17'd63782;
    value[5038] = 17'd63769;
    value[5039] = 17'd63755;
    value[5040] = 17'd63742;
    value[5041] = 17'd63728;
    value[5042] = 17'd63715;
    value[5043] = 17'd63702;
    value[5044] = 17'd63688;
    value[5045] = 17'd63675;
    value[5046] = 17'd63661;
    value[5047] = 17'd63648;
    value[5048] = 17'd63634;
    value[5049] = 17'd63621;
    value[5050] = 17'd63607;
    value[5051] = 17'd63594;
    value[5052] = 17'd63580;
    value[5053] = 17'd63567;
    value[5054] = 17'd63553;
    value[5055] = 17'd63540;
    value[5056] = 17'd63526;
    value[5057] = 17'd63513;
    value[5058] = 17'd63500;
    value[5059] = 17'd63486;
    value[5060] = 17'd63473;
    value[5061] = 17'd63459;
    value[5062] = 17'd63446;
    value[5063] = 17'd63432;
    value[5064] = 17'd63419;
    value[5065] = 17'd63405;
    value[5066] = 17'd63392;
    value[5067] = 17'd63378;
    value[5068] = 17'd63365;
    value[5069] = 17'd63351;
    value[5070] = 17'd63338;
    value[5071] = 17'd63324;
    value[5072] = 17'd63311;
    value[5073] = 17'd63297;
    value[5074] = 17'd63284;
    value[5075] = 17'd63270;
    value[5076] = 17'd63257;
    value[5077] = 17'd63243;
    value[5078] = 17'd63229;
    value[5079] = 17'd63216;
    value[5080] = 17'd63202;
    value[5081] = 17'd63189;
    value[5082] = 17'd63175;
    value[5083] = 17'd63162;
    value[5084] = 17'd63148;
    value[5085] = 17'd63135;
    value[5086] = 17'd63121;
    value[5087] = 17'd63108;
    value[5088] = 17'd63094;
    value[5089] = 17'd63081;
    value[5090] = 17'd63067;
    value[5091] = 17'd63054;
    value[5092] = 17'd63040;
    value[5093] = 17'd63026;
    value[5094] = 17'd63013;
    value[5095] = 17'd62999;
    value[5096] = 17'd62986;
    value[5097] = 17'd62972;
    value[5098] = 17'd62959;
    value[5099] = 17'd62945;
    value[5100] = 17'd62932;
    value[5101] = 17'd62918;
    value[5102] = 17'd62904;
    value[5103] = 17'd62891;
    value[5104] = 17'd62877;
    value[5105] = 17'd62864;
    value[5106] = 17'd62850;
    value[5107] = 17'd62837;
    value[5108] = 17'd62823;
    value[5109] = 17'd62809;
    value[5110] = 17'd62796;
    value[5111] = 17'd62782;
    value[5112] = 17'd62769;
    value[5113] = 17'd62755;
    value[5114] = 17'd62741;
    value[5115] = 17'd62728;
    value[5116] = 17'd62714;
    value[5117] = 17'd62701;
    value[5118] = 17'd62687;
    value[5119] = 17'd62673;
    value[5120] = 17'd62660;
    value[5121] = 17'd62646;
    value[5122] = 17'd62633;
    value[5123] = 17'd62619;
    value[5124] = 17'd62605;
    value[5125] = 17'd62592;
    value[5126] = 17'd62578;
    value[5127] = 17'd62565;
    value[5128] = 17'd62551;
    value[5129] = 17'd62537;
    value[5130] = 17'd62524;
    value[5131] = 17'd62510;
    value[5132] = 17'd62497;
    value[5133] = 17'd62483;
    value[5134] = 17'd62469;
    value[5135] = 17'd62456;
    value[5136] = 17'd62442;
    value[5137] = 17'd62428;
    value[5138] = 17'd62415;
    value[5139] = 17'd62401;
    value[5140] = 17'd62387;
    value[5141] = 17'd62374;
    value[5142] = 17'd62360;
    value[5143] = 17'd62347;
    value[5144] = 17'd62333;
    value[5145] = 17'd62319;
    value[5146] = 17'd62306;
    value[5147] = 17'd62292;
    value[5148] = 17'd62278;
    value[5149] = 17'd62265;
    value[5150] = 17'd62251;
    value[5151] = 17'd62237;
    value[5152] = 17'd62224;
    value[5153] = 17'd62210;
    value[5154] = 17'd62196;
    value[5155] = 17'd62183;
    value[5156] = 17'd62169;
    value[5157] = 17'd62155;
    value[5158] = 17'd62142;
    value[5159] = 17'd62128;
    value[5160] = 17'd62114;
    value[5161] = 17'd62101;
    value[5162] = 17'd62087;
    value[5163] = 17'd62073;
    value[5164] = 17'd62060;
    value[5165] = 17'd62046;
    value[5166] = 17'd62032;
    value[5167] = 17'd62018;
    value[5168] = 17'd62005;
    value[5169] = 17'd61991;
    value[5170] = 17'd61977;
    value[5171] = 17'd61964;
    value[5172] = 17'd61950;
    value[5173] = 17'd61936;
    value[5174] = 17'd61923;
    value[5175] = 17'd61909;
    value[5176] = 17'd61895;
    value[5177] = 17'd61881;
    value[5178] = 17'd61868;
    value[5179] = 17'd61854;
    value[5180] = 17'd61840;
    value[5181] = 17'd61827;
    value[5182] = 17'd61813;
    value[5183] = 17'd61799;
    value[5184] = 17'd61785;
    value[5185] = 17'd61772;
    value[5186] = 17'd61758;
    value[5187] = 17'd61744;
    value[5188] = 17'd61731;
    value[5189] = 17'd61717;
    value[5190] = 17'd61703;
    value[5191] = 17'd61689;
    value[5192] = 17'd61676;
    value[5193] = 17'd61662;
    value[5194] = 17'd61648;
    value[5195] = 17'd61634;
    value[5196] = 17'd61621;
    value[5197] = 17'd61607;
    value[5198] = 17'd61593;
    value[5199] = 17'd61579;
    value[5200] = 17'd61566;
    value[5201] = 17'd61552;
    value[5202] = 17'd61538;
    value[5203] = 17'd61524;
    value[5204] = 17'd61511;
    value[5205] = 17'd61497;
    value[5206] = 17'd61483;
    value[5207] = 17'd61469;
    value[5208] = 17'd61456;
    value[5209] = 17'd61442;
    value[5210] = 17'd61428;
    value[5211] = 17'd61414;
    value[5212] = 17'd61400;
    value[5213] = 17'd61387;
    value[5214] = 17'd61373;
    value[5215] = 17'd61359;
    value[5216] = 17'd61345;
    value[5217] = 17'd61332;
    value[5218] = 17'd61318;
    value[5219] = 17'd61304;
    value[5220] = 17'd61290;
    value[5221] = 17'd61276;
    value[5222] = 17'd61263;
    value[5223] = 17'd61249;
    value[5224] = 17'd61235;
    value[5225] = 17'd61221;
    value[5226] = 17'd61207;
    value[5227] = 17'd61194;
    value[5228] = 17'd61180;
    value[5229] = 17'd61166;
    value[5230] = 17'd61152;
    value[5231] = 17'd61138;
    value[5232] = 17'd61125;
    value[5233] = 17'd61111;
    value[5234] = 17'd61097;
    value[5235] = 17'd61083;
    value[5236] = 17'd61069;
    value[5237] = 17'd61055;
    value[5238] = 17'd61042;
    value[5239] = 17'd61028;
    value[5240] = 17'd61014;
    value[5241] = 17'd61000;
    value[5242] = 17'd60986;
    value[5243] = 17'd60973;
    value[5244] = 17'd60959;
    value[5245] = 17'd60945;
    value[5246] = 17'd60931;
    value[5247] = 17'd60917;
    value[5248] = 17'd60903;
    value[5249] = 17'd60889;
    value[5250] = 17'd60876;
    value[5251] = 17'd60862;
    value[5252] = 17'd60848;
    value[5253] = 17'd60834;
    value[5254] = 17'd60820;
    value[5255] = 17'd60806;
    value[5256] = 17'd60793;
    value[5257] = 17'd60779;
    value[5258] = 17'd60765;
    value[5259] = 17'd60751;
    value[5260] = 17'd60737;
    value[5261] = 17'd60723;
    value[5262] = 17'd60709;
    value[5263] = 17'd60695;
    value[5264] = 17'd60682;
    value[5265] = 17'd60668;
    value[5266] = 17'd60654;
    value[5267] = 17'd60640;
    value[5268] = 17'd60626;
    value[5269] = 17'd60612;
    value[5270] = 17'd60598;
    value[5271] = 17'd60584;
    value[5272] = 17'd60571;
    value[5273] = 17'd60557;
    value[5274] = 17'd60543;
    value[5275] = 17'd60529;
    value[5276] = 17'd60515;
    value[5277] = 17'd60501;
    value[5278] = 17'd60487;
    value[5279] = 17'd60473;
    value[5280] = 17'd60459;
    value[5281] = 17'd60446;
    value[5282] = 17'd60432;
    value[5283] = 17'd60418;
    value[5284] = 17'd60404;
    value[5285] = 17'd60390;
    value[5286] = 17'd60376;
    value[5287] = 17'd60362;
    value[5288] = 17'd60348;
    value[5289] = 17'd60334;
    value[5290] = 17'd60320;
    value[5291] = 17'd60306;
    value[5292] = 17'd60292;
    value[5293] = 17'd60279;
    value[5294] = 17'd60265;
    value[5295] = 17'd60251;
    value[5296] = 17'd60237;
    value[5297] = 17'd60223;
    value[5298] = 17'd60209;
    value[5299] = 17'd60195;
    value[5300] = 17'd60181;
    value[5301] = 17'd60167;
    value[5302] = 17'd60153;
    value[5303] = 17'd60139;
    value[5304] = 17'd60125;
    value[5305] = 17'd60111;
    value[5306] = 17'd60097;
    value[5307] = 17'd60083;
    value[5308] = 17'd60069;
    value[5309] = 17'd60055;
    value[5310] = 17'd60042;
    value[5311] = 17'd60028;
    value[5312] = 17'd60014;
    value[5313] = 17'd60000;
    value[5314] = 17'd59986;
    value[5315] = 17'd59972;
    value[5316] = 17'd59958;
    value[5317] = 17'd59944;
    value[5318] = 17'd59930;
    value[5319] = 17'd59916;
    value[5320] = 17'd59902;
    value[5321] = 17'd59888;
    value[5322] = 17'd59874;
    value[5323] = 17'd59860;
    value[5324] = 17'd59846;
    value[5325] = 17'd59832;
    value[5326] = 17'd59818;
    value[5327] = 17'd59804;
    value[5328] = 17'd59790;
    value[5329] = 17'd59776;
    value[5330] = 17'd59762;
    value[5331] = 17'd59748;
    value[5332] = 17'd59734;
    value[5333] = 17'd59720;
    value[5334] = 17'd59706;
    value[5335] = 17'd59692;
    value[5336] = 17'd59678;
    value[5337] = 17'd59664;
    value[5338] = 17'd59650;
    value[5339] = 17'd59636;
    value[5340] = 17'd59622;
    value[5341] = 17'd59608;
    value[5342] = 17'd59594;
    value[5343] = 17'd59580;
    value[5344] = 17'd59566;
    value[5345] = 17'd59552;
    value[5346] = 17'd59538;
    value[5347] = 17'd59524;
    value[5348] = 17'd59510;
    value[5349] = 17'd59496;
    value[5350] = 17'd59482;
    value[5351] = 17'd59468;
    value[5352] = 17'd59454;
    value[5353] = 17'd59440;
    value[5354] = 17'd59426;
    value[5355] = 17'd59412;
    value[5356] = 17'd59398;
    value[5357] = 17'd59384;
    value[5358] = 17'd59369;
    value[5359] = 17'd59355;
    value[5360] = 17'd59341;
    value[5361] = 17'd59327;
    value[5362] = 17'd59313;
    value[5363] = 17'd59299;
    value[5364] = 17'd59285;
    value[5365] = 17'd59271;
    value[5366] = 17'd59257;
    value[5367] = 17'd59243;
    value[5368] = 17'd59229;
    value[5369] = 17'd59215;
    value[5370] = 17'd59201;
    value[5371] = 17'd59187;
    value[5372] = 17'd59173;
    value[5373] = 17'd59159;
    value[5374] = 17'd59145;
    value[5375] = 17'd59130;
    value[5376] = 17'd59116;
    value[5377] = 17'd59102;
    value[5378] = 17'd59088;
    value[5379] = 17'd59074;
    value[5380] = 17'd59060;
    value[5381] = 17'd59046;
    value[5382] = 17'd59032;
    value[5383] = 17'd59018;
    value[5384] = 17'd59004;
    value[5385] = 17'd58990;
    value[5386] = 17'd58976;
    value[5387] = 17'd58961;
    value[5388] = 17'd58947;
    value[5389] = 17'd58933;
    value[5390] = 17'd58919;
    value[5391] = 17'd58905;
    value[5392] = 17'd58891;
    value[5393] = 17'd58877;
    value[5394] = 17'd58863;
    value[5395] = 17'd58849;
    value[5396] = 17'd58834;
    value[5397] = 17'd58820;
    value[5398] = 17'd58806;
    value[5399] = 17'd58792;
    value[5400] = 17'd58778;
    value[5401] = 17'd58764;
    value[5402] = 17'd58750;
    value[5403] = 17'd58736;
    value[5404] = 17'd58722;
    value[5405] = 17'd58707;
    value[5406] = 17'd58693;
    value[5407] = 17'd58679;
    value[5408] = 17'd58665;
    value[5409] = 17'd58651;
    value[5410] = 17'd58637;
    value[5411] = 17'd58623;
    value[5412] = 17'd58608;
    value[5413] = 17'd58594;
    value[5414] = 17'd58580;
    value[5415] = 17'd58566;
    value[5416] = 17'd58552;
    value[5417] = 17'd58538;
    value[5418] = 17'd58524;
    value[5419] = 17'd58509;
    value[5420] = 17'd58495;
    value[5421] = 17'd58481;
    value[5422] = 17'd58467;
    value[5423] = 17'd58453;
    value[5424] = 17'd58439;
    value[5425] = 17'd58424;
    value[5426] = 17'd58410;
    value[5427] = 17'd58396;
    value[5428] = 17'd58382;
    value[5429] = 17'd58368;
    value[5430] = 17'd58354;
    value[5431] = 17'd58339;
    value[5432] = 17'd58325;
    value[5433] = 17'd58311;
    value[5434] = 17'd58297;
    value[5435] = 17'd58283;
    value[5436] = 17'd58269;
    value[5437] = 17'd58254;
    value[5438] = 17'd58240;
    value[5439] = 17'd58226;
    value[5440] = 17'd58212;
    value[5441] = 17'd58198;
    value[5442] = 17'd58183;
    value[5443] = 17'd58169;
    value[5444] = 17'd58155;
    value[5445] = 17'd58141;
    value[5446] = 17'd58127;
    value[5447] = 17'd58112;
    value[5448] = 17'd58098;
    value[5449] = 17'd58084;
    value[5450] = 17'd58070;
    value[5451] = 17'd58056;
    value[5452] = 17'd58041;
    value[5453] = 17'd58027;
    value[5454] = 17'd58013;
    value[5455] = 17'd57999;
    value[5456] = 17'd57985;
    value[5457] = 17'd57970;
    value[5458] = 17'd57956;
    value[5459] = 17'd57942;
    value[5460] = 17'd57928;
    value[5461] = 17'd57913;
    value[5462] = 17'd57899;
    value[5463] = 17'd57885;
    value[5464] = 17'd57871;
    value[5465] = 17'd57856;
    value[5466] = 17'd57842;
    value[5467] = 17'd57828;
    value[5468] = 17'd57814;
    value[5469] = 17'd57800;
    value[5470] = 17'd57785;
    value[5471] = 17'd57771;
    value[5472] = 17'd57757;
    value[5473] = 17'd57743;
    value[5474] = 17'd57728;
    value[5475] = 17'd57714;
    value[5476] = 17'd57700;
    value[5477] = 17'd57686;
    value[5478] = 17'd57671;
    value[5479] = 17'd57657;
    value[5480] = 17'd57643;
    value[5481] = 17'd57628;
    value[5482] = 17'd57614;
    value[5483] = 17'd57600;
    value[5484] = 17'd57586;
    value[5485] = 17'd57571;
    value[5486] = 17'd57557;
    value[5487] = 17'd57543;
    value[5488] = 17'd57529;
    value[5489] = 17'd57514;
    value[5490] = 17'd57500;
    value[5491] = 17'd57486;
    value[5492] = 17'd57471;
    value[5493] = 17'd57457;
    value[5494] = 17'd57443;
    value[5495] = 17'd57429;
    value[5496] = 17'd57414;
    value[5497] = 17'd57400;
    value[5498] = 17'd57386;
    value[5499] = 17'd57371;
    value[5500] = 17'd57357;
    value[5501] = 17'd57343;
    value[5502] = 17'd57329;
    value[5503] = 17'd57314;
    value[5504] = 17'd57300;
    value[5505] = 17'd57286;
    value[5506] = 17'd57271;
    value[5507] = 17'd57257;
    value[5508] = 17'd57243;
    value[5509] = 17'd57228;
    value[5510] = 17'd57214;
    value[5511] = 17'd57200;
    value[5512] = 17'd57185;
    value[5513] = 17'd57171;
    value[5514] = 17'd57157;
    value[5515] = 17'd57142;
    value[5516] = 17'd57128;
    value[5517] = 17'd57114;
    value[5518] = 17'd57100;
    value[5519] = 17'd57085;
    value[5520] = 17'd57071;
    value[5521] = 17'd57057;
    value[5522] = 17'd57042;
    value[5523] = 17'd57028;
    value[5524] = 17'd57014;
    value[5525] = 17'd56999;
    value[5526] = 17'd56985;
    value[5527] = 17'd56970;
    value[5528] = 17'd56956;
    value[5529] = 17'd56942;
    value[5530] = 17'd56927;
    value[5531] = 17'd56913;
    value[5532] = 17'd56899;
    value[5533] = 17'd56884;
    value[5534] = 17'd56870;
    value[5535] = 17'd56856;
    value[5536] = 17'd56841;
    value[5537] = 17'd56827;
    value[5538] = 17'd56813;
    value[5539] = 17'd56798;
    value[5540] = 17'd56784;
    value[5541] = 17'd56770;
    value[5542] = 17'd56755;
    value[5543] = 17'd56741;
    value[5544] = 17'd56726;
    value[5545] = 17'd56712;
    value[5546] = 17'd56698;
    value[5547] = 17'd56683;
    value[5548] = 17'd56669;
    value[5549] = 17'd56655;
    value[5550] = 17'd56640;
    value[5551] = 17'd56626;
    value[5552] = 17'd56611;
    value[5553] = 17'd56597;
    value[5554] = 17'd56583;
    value[5555] = 17'd56568;
    value[5556] = 17'd56554;
    value[5557] = 17'd56539;
    value[5558] = 17'd56525;
    value[5559] = 17'd56511;
    value[5560] = 17'd56496;
    value[5561] = 17'd56482;
    value[5562] = 17'd56467;
    value[5563] = 17'd56453;
    value[5564] = 17'd56439;
    value[5565] = 17'd56424;
    value[5566] = 17'd56410;
    value[5567] = 17'd56395;
    value[5568] = 17'd56381;
    value[5569] = 17'd56367;
    value[5570] = 17'd56352;
    value[5571] = 17'd56338;
    value[5572] = 17'd56323;
    value[5573] = 17'd56309;
    value[5574] = 17'd56294;
    value[5575] = 17'd56280;
    value[5576] = 17'd56266;
    value[5577] = 17'd56251;
    value[5578] = 17'd56237;
    value[5579] = 17'd56222;
    value[5580] = 17'd56208;
    value[5581] = 17'd56193;
    value[5582] = 17'd56179;
    value[5583] = 17'd56165;
    value[5584] = 17'd56150;
    value[5585] = 17'd56136;
    value[5586] = 17'd56121;
    value[5587] = 17'd56107;
    value[5588] = 17'd56092;
    value[5589] = 17'd56078;
    value[5590] = 17'd56063;
    value[5591] = 17'd56049;
    value[5592] = 17'd56034;
    value[5593] = 17'd56020;
    value[5594] = 17'd56006;
    value[5595] = 17'd55991;
    value[5596] = 17'd55977;
    value[5597] = 17'd55962;
    value[5598] = 17'd55948;
    value[5599] = 17'd55933;
    value[5600] = 17'd55919;
    value[5601] = 17'd55904;
    value[5602] = 17'd55890;
    value[5603] = 17'd55875;
    value[5604] = 17'd55861;
    value[5605] = 17'd55846;
    value[5606] = 17'd55832;
    value[5607] = 17'd55817;
    value[5608] = 17'd55803;
    value[5609] = 17'd55788;
    value[5610] = 17'd55774;
    value[5611] = 17'd55760;
    value[5612] = 17'd55745;
    value[5613] = 17'd55731;
    value[5614] = 17'd55716;
    value[5615] = 17'd55702;
    value[5616] = 17'd55687;
    value[5617] = 17'd55673;
    value[5618] = 17'd55658;
    value[5619] = 17'd55644;
    value[5620] = 17'd55629;
    value[5621] = 17'd55615;
    value[5622] = 17'd55600;
    value[5623] = 17'd55586;
    value[5624] = 17'd55571;
    value[5625] = 17'd55557;
    value[5626] = 17'd55542;
    value[5627] = 17'd55527;
    value[5628] = 17'd55513;
    value[5629] = 17'd55498;
    value[5630] = 17'd55484;
    value[5631] = 17'd55469;
    value[5632] = 17'd55455;
    value[5633] = 17'd55440;
    value[5634] = 17'd55426;
    value[5635] = 17'd55411;
    value[5636] = 17'd55397;
    value[5637] = 17'd55382;
    value[5638] = 17'd55368;
    value[5639] = 17'd55353;
    value[5640] = 17'd55339;
    value[5641] = 17'd55324;
    value[5642] = 17'd55310;
    value[5643] = 17'd55295;
    value[5644] = 17'd55280;
    value[5645] = 17'd55266;
    value[5646] = 17'd55251;
    value[5647] = 17'd55237;
    value[5648] = 17'd55222;
    value[5649] = 17'd55208;
    value[5650] = 17'd55193;
    value[5651] = 17'd55179;
    value[5652] = 17'd55164;
    value[5653] = 17'd55150;
    value[5654] = 17'd55135;
    value[5655] = 17'd55120;
    value[5656] = 17'd55106;
    value[5657] = 17'd55091;
    value[5658] = 17'd55077;
    value[5659] = 17'd55062;
    value[5660] = 17'd55048;
    value[5661] = 17'd55033;
    value[5662] = 17'd55018;
    value[5663] = 17'd55004;
    value[5664] = 17'd54989;
    value[5665] = 17'd54975;
    value[5666] = 17'd54960;
    value[5667] = 17'd54946;
    value[5668] = 17'd54931;
    value[5669] = 17'd54916;
    value[5670] = 17'd54902;
    value[5671] = 17'd54887;
    value[5672] = 17'd54873;
    value[5673] = 17'd54858;
    value[5674] = 17'd54843;
    value[5675] = 17'd54829;
    value[5676] = 17'd54814;
    value[5677] = 17'd54800;
    value[5678] = 17'd54785;
    value[5679] = 17'd54770;
    value[5680] = 17'd54756;
    value[5681] = 17'd54741;
    value[5682] = 17'd54727;
    value[5683] = 17'd54712;
    value[5684] = 17'd54697;
    value[5685] = 17'd54683;
    value[5686] = 17'd54668;
    value[5687] = 17'd54654;
    value[5688] = 17'd54639;
    value[5689] = 17'd54624;
    value[5690] = 17'd54610;
    value[5691] = 17'd54595;
    value[5692] = 17'd54580;
    value[5693] = 17'd54566;
    value[5694] = 17'd54551;
    value[5695] = 17'd54537;
    value[5696] = 17'd54522;
    value[5697] = 17'd54507;
    value[5698] = 17'd54493;
    value[5699] = 17'd54478;
    value[5700] = 17'd54463;
    value[5701] = 17'd54449;
    value[5702] = 17'd54434;
    value[5703] = 17'd54419;
    value[5704] = 17'd54405;
    value[5705] = 17'd54390;
    value[5706] = 17'd54376;
    value[5707] = 17'd54361;
    value[5708] = 17'd54346;
    value[5709] = 17'd54332;
    value[5710] = 17'd54317;
    value[5711] = 17'd54302;
    value[5712] = 17'd54288;
    value[5713] = 17'd54273;
    value[5714] = 17'd54258;
    value[5715] = 17'd54244;
    value[5716] = 17'd54229;
    value[5717] = 17'd54214;
    value[5718] = 17'd54200;
    value[5719] = 17'd54185;
    value[5720] = 17'd54170;
    value[5721] = 17'd54156;
    value[5722] = 17'd54141;
    value[5723] = 17'd54126;
    value[5724] = 17'd54112;
    value[5725] = 17'd54097;
    value[5726] = 17'd54082;
    value[5727] = 17'd54068;
    value[5728] = 17'd54053;
    value[5729] = 17'd54038;
    value[5730] = 17'd54024;
    value[5731] = 17'd54009;
    value[5732] = 17'd53994;
    value[5733] = 17'd53979;
    value[5734] = 17'd53965;
    value[5735] = 17'd53950;
    value[5736] = 17'd53935;
    value[5737] = 17'd53921;
    value[5738] = 17'd53906;
    value[5739] = 17'd53891;
    value[5740] = 17'd53877;
    value[5741] = 17'd53862;
    value[5742] = 17'd53847;
    value[5743] = 17'd53832;
    value[5744] = 17'd53818;
    value[5745] = 17'd53803;
    value[5746] = 17'd53788;
    value[5747] = 17'd53774;
    value[5748] = 17'd53759;
    value[5749] = 17'd53744;
    value[5750] = 17'd53729;
    value[5751] = 17'd53715;
    value[5752] = 17'd53700;
    value[5753] = 17'd53685;
    value[5754] = 17'd53671;
    value[5755] = 17'd53656;
    value[5756] = 17'd53641;
    value[5757] = 17'd53626;
    value[5758] = 17'd53612;
    value[5759] = 17'd53597;
    value[5760] = 17'd53582;
    value[5761] = 17'd53567;
    value[5762] = 17'd53553;
    value[5763] = 17'd53538;
    value[5764] = 17'd53523;
    value[5765] = 17'd53508;
    value[5766] = 17'd53494;
    value[5767] = 17'd53479;
    value[5768] = 17'd53464;
    value[5769] = 17'd53449;
    value[5770] = 17'd53435;
    value[5771] = 17'd53420;
    value[5772] = 17'd53405;
    value[5773] = 17'd53390;
    value[5774] = 17'd53376;
    value[5775] = 17'd53361;
    value[5776] = 17'd53346;
    value[5777] = 17'd53331;
    value[5778] = 17'd53317;
    value[5779] = 17'd53302;
    value[5780] = 17'd53287;
    value[5781] = 17'd53272;
    value[5782] = 17'd53258;
    value[5783] = 17'd53243;
    value[5784] = 17'd53228;
    value[5785] = 17'd53213;
    value[5786] = 17'd53198;
    value[5787] = 17'd53184;
    value[5788] = 17'd53169;
    value[5789] = 17'd53154;
    value[5790] = 17'd53139;
    value[5791] = 17'd53125;
    value[5792] = 17'd53110;
    value[5793] = 17'd53095;
    value[5794] = 17'd53080;
    value[5795] = 17'd53065;
    value[5796] = 17'd53051;
    value[5797] = 17'd53036;
    value[5798] = 17'd53021;
    value[5799] = 17'd53006;
    value[5800] = 17'd52991;
    value[5801] = 17'd52977;
    value[5802] = 17'd52962;
    value[5803] = 17'd52947;
    value[5804] = 17'd52932;
    value[5805] = 17'd52917;
    value[5806] = 17'd52903;
    value[5807] = 17'd52888;
    value[5808] = 17'd52873;
    value[5809] = 17'd52858;
    value[5810] = 17'd52843;
    value[5811] = 17'd52829;
    value[5812] = 17'd52814;
    value[5813] = 17'd52799;
    value[5814] = 17'd52784;
    value[5815] = 17'd52769;
    value[5816] = 17'd52754;
    value[5817] = 17'd52740;
    value[5818] = 17'd52725;
    value[5819] = 17'd52710;
    value[5820] = 17'd52695;
    value[5821] = 17'd52680;
    value[5822] = 17'd52665;
    value[5823] = 17'd52651;
    value[5824] = 17'd52636;
    value[5825] = 17'd52621;
    value[5826] = 17'd52606;
    value[5827] = 17'd52591;
    value[5828] = 17'd52576;
    value[5829] = 17'd52562;
    value[5830] = 17'd52547;
    value[5831] = 17'd52532;
    value[5832] = 17'd52517;
    value[5833] = 17'd52502;
    value[5834] = 17'd52487;
    value[5835] = 17'd52472;
    value[5836] = 17'd52458;
    value[5837] = 17'd52443;
    value[5838] = 17'd52428;
    value[5839] = 17'd52413;
    value[5840] = 17'd52398;
    value[5841] = 17'd52383;
    value[5842] = 17'd52368;
    value[5843] = 17'd52353;
    value[5844] = 17'd52339;
    value[5845] = 17'd52324;
    value[5846] = 17'd52309;
    value[5847] = 17'd52294;
    value[5848] = 17'd52279;
    value[5849] = 17'd52264;
    value[5850] = 17'd52249;
    value[5851] = 17'd52234;
    value[5852] = 17'd52220;
    value[5853] = 17'd52205;
    value[5854] = 17'd52190;
    value[5855] = 17'd52175;
    value[5856] = 17'd52160;
    value[5857] = 17'd52145;
    value[5858] = 17'd52130;
    value[5859] = 17'd52115;
    value[5860] = 17'd52100;
    value[5861] = 17'd52086;
    value[5862] = 17'd52071;
    value[5863] = 17'd52056;
    value[5864] = 17'd52041;
    value[5865] = 17'd52026;
    value[5866] = 17'd52011;
    value[5867] = 17'd51996;
    value[5868] = 17'd51981;
    value[5869] = 17'd51966;
    value[5870] = 17'd51951;
    value[5871] = 17'd51936;
    value[5872] = 17'd51922;
    value[5873] = 17'd51907;
    value[5874] = 17'd51892;
    value[5875] = 17'd51877;
    value[5876] = 17'd51862;
    value[5877] = 17'd51847;
    value[5878] = 17'd51832;
    value[5879] = 17'd51817;
    value[5880] = 17'd51802;
    value[5881] = 17'd51787;
    value[5882] = 17'd51772;
    value[5883] = 17'd51757;
    value[5884] = 17'd51742;
    value[5885] = 17'd51728;
    value[5886] = 17'd51713;
    value[5887] = 17'd51698;
    value[5888] = 17'd51683;
    value[5889] = 17'd51668;
    value[5890] = 17'd51653;
    value[5891] = 17'd51638;
    value[5892] = 17'd51623;
    value[5893] = 17'd51608;
    value[5894] = 17'd51593;
    value[5895] = 17'd51578;
    value[5896] = 17'd51563;
    value[5897] = 17'd51548;
    value[5898] = 17'd51533;
    value[5899] = 17'd51518;
    value[5900] = 17'd51503;
    value[5901] = 17'd51488;
    value[5902] = 17'd51473;
    value[5903] = 17'd51458;
    value[5904] = 17'd51443;
    value[5905] = 17'd51428;
    value[5906] = 17'd51414;
    value[5907] = 17'd51399;
    value[5908] = 17'd51384;
    value[5909] = 17'd51369;
    value[5910] = 17'd51354;
    value[5911] = 17'd51339;
    value[5912] = 17'd51324;
    value[5913] = 17'd51309;
    value[5914] = 17'd51294;
    value[5915] = 17'd51279;
    value[5916] = 17'd51264;
    value[5917] = 17'd51249;
    value[5918] = 17'd51234;
    value[5919] = 17'd51219;
    value[5920] = 17'd51204;
    value[5921] = 17'd51189;
    value[5922] = 17'd51174;
    value[5923] = 17'd51159;
    value[5924] = 17'd51144;
    value[5925] = 17'd51129;
    value[5926] = 17'd51114;
    value[5927] = 17'd51099;
    value[5928] = 17'd51084;
    value[5929] = 17'd51069;
    value[5930] = 17'd51054;
    value[5931] = 17'd51039;
    value[5932] = 17'd51024;
    value[5933] = 17'd51009;
    value[5934] = 17'd50994;
    value[5935] = 17'd50979;
    value[5936] = 17'd50964;
    value[5937] = 17'd50949;
    value[5938] = 17'd50934;
    value[5939] = 17'd50919;
    value[5940] = 17'd50904;
    value[5941] = 17'd50889;
    value[5942] = 17'd50874;
    value[5943] = 17'd50859;
    value[5944] = 17'd50844;
    value[5945] = 17'd50829;
    value[5946] = 17'd50813;
    value[5947] = 17'd50798;
    value[5948] = 17'd50783;
    value[5949] = 17'd50768;
    value[5950] = 17'd50753;
    value[5951] = 17'd50738;
    value[5952] = 17'd50723;
    value[5953] = 17'd50708;
    value[5954] = 17'd50693;
    value[5955] = 17'd50678;
    value[5956] = 17'd50663;
    value[5957] = 17'd50648;
    value[5958] = 17'd50633;
    value[5959] = 17'd50618;
    value[5960] = 17'd50603;
    value[5961] = 17'd50588;
    value[5962] = 17'd50573;
    value[5963] = 17'd50558;
    value[5964] = 17'd50543;
    value[5965] = 17'd50528;
    value[5966] = 17'd50513;
    value[5967] = 17'd50497;
    value[5968] = 17'd50482;
    value[5969] = 17'd50467;
    value[5970] = 17'd50452;
    value[5971] = 17'd50437;
    value[5972] = 17'd50422;
    value[5973] = 17'd50407;
    value[5974] = 17'd50392;
    value[5975] = 17'd50377;
    value[5976] = 17'd50362;
    value[5977] = 17'd50347;
    value[5978] = 17'd50332;
    value[5979] = 17'd50317;
    value[5980] = 17'd50301;
    value[5981] = 17'd50286;
    value[5982] = 17'd50271;
    value[5983] = 17'd50256;
    value[5984] = 17'd50241;
    value[5985] = 17'd50226;
    value[5986] = 17'd50211;
    value[5987] = 17'd50196;
    value[5988] = 17'd50181;
    value[5989] = 17'd50166;
    value[5990] = 17'd50151;
    value[5991] = 17'd50135;
    value[5992] = 17'd50120;
    value[5993] = 17'd50105;
    value[5994] = 17'd50090;
    value[5995] = 17'd50075;
    value[5996] = 17'd50060;
    value[5997] = 17'd50045;
    value[5998] = 17'd50030;
    value[5999] = 17'd50015;
    value[6000] = 17'd50000;
    value[6001] = 17'd49984;
    value[6002] = 17'd49969;
    value[6003] = 17'd49954;
    value[6004] = 17'd49939;
    value[6005] = 17'd49924;
    value[6006] = 17'd49909;
    value[6007] = 17'd49894;
    value[6008] = 17'd49879;
    value[6009] = 17'd49863;
    value[6010] = 17'd49848;
    value[6011] = 17'd49833;
    value[6012] = 17'd49818;
    value[6013] = 17'd49803;
    value[6014] = 17'd49788;
    value[6015] = 17'd49773;
    value[6016] = 17'd49757;
    value[6017] = 17'd49742;
    value[6018] = 17'd49727;
    value[6019] = 17'd49712;
    value[6020] = 17'd49697;
    value[6021] = 17'd49682;
    value[6022] = 17'd49667;
    value[6023] = 17'd49651;
    value[6024] = 17'd49636;
    value[6025] = 17'd49621;
    value[6026] = 17'd49606;
    value[6027] = 17'd49591;
    value[6028] = 17'd49576;
    value[6029] = 17'd49561;
    value[6030] = 17'd49545;
    value[6031] = 17'd49530;
    value[6032] = 17'd49515;
    value[6033] = 17'd49500;
    value[6034] = 17'd49485;
    value[6035] = 17'd49470;
    value[6036] = 17'd49454;
    value[6037] = 17'd49439;
    value[6038] = 17'd49424;
    value[6039] = 17'd49409;
    value[6040] = 17'd49394;
    value[6041] = 17'd49379;
    value[6042] = 17'd49363;
    value[6043] = 17'd49348;
    value[6044] = 17'd49333;
    value[6045] = 17'd49318;
    value[6046] = 17'd49303;
    value[6047] = 17'd49287;
    value[6048] = 17'd49272;
    value[6049] = 17'd49257;
    value[6050] = 17'd49242;
    value[6051] = 17'd49227;
    value[6052] = 17'd49211;
    value[6053] = 17'd49196;
    value[6054] = 17'd49181;
    value[6055] = 17'd49166;
    value[6056] = 17'd49151;
    value[6057] = 17'd49135;
    value[6058] = 17'd49120;
    value[6059] = 17'd49105;
    value[6060] = 17'd49090;
    value[6061] = 17'd49075;
    value[6062] = 17'd49059;
    value[6063] = 17'd49044;
    value[6064] = 17'd49029;
    value[6065] = 17'd49014;
    value[6066] = 17'd48999;
    value[6067] = 17'd48983;
    value[6068] = 17'd48968;
    value[6069] = 17'd48953;
    value[6070] = 17'd48938;
    value[6071] = 17'd48923;
    value[6072] = 17'd48907;
    value[6073] = 17'd48892;
    value[6074] = 17'd48877;
    value[6075] = 17'd48862;
    value[6076] = 17'd48846;
    value[6077] = 17'd48831;
    value[6078] = 17'd48816;
    value[6079] = 17'd48801;
    value[6080] = 17'd48785;
    value[6081] = 17'd48770;
    value[6082] = 17'd48755;
    value[6083] = 17'd48740;
    value[6084] = 17'd48725;
    value[6085] = 17'd48709;
    value[6086] = 17'd48694;
    value[6087] = 17'd48679;
    value[6088] = 17'd48664;
    value[6089] = 17'd48648;
    value[6090] = 17'd48633;
    value[6091] = 17'd48618;
    value[6092] = 17'd48603;
    value[6093] = 17'd48587;
    value[6094] = 17'd48572;
    value[6095] = 17'd48557;
    value[6096] = 17'd48542;
    value[6097] = 17'd48526;
    value[6098] = 17'd48511;
    value[6099] = 17'd48496;
    value[6100] = 17'd48480;
    value[6101] = 17'd48465;
    value[6102] = 17'd48450;
    value[6103] = 17'd48435;
    value[6104] = 17'd48419;
    value[6105] = 17'd48404;
    value[6106] = 17'd48389;
    value[6107] = 17'd48374;
    value[6108] = 17'd48358;
    value[6109] = 17'd48343;
    value[6110] = 17'd48328;
    value[6111] = 17'd48312;
    value[6112] = 17'd48297;
    value[6113] = 17'd48282;
    value[6114] = 17'd48267;
    value[6115] = 17'd48251;
    value[6116] = 17'd48236;
    value[6117] = 17'd48221;
    value[6118] = 17'd48205;
    value[6119] = 17'd48190;
    value[6120] = 17'd48175;
    value[6121] = 17'd48160;
    value[6122] = 17'd48144;
    value[6123] = 17'd48129;
    value[6124] = 17'd48114;
    value[6125] = 17'd48098;
    value[6126] = 17'd48083;
    value[6127] = 17'd48068;
    value[6128] = 17'd48052;
    value[6129] = 17'd48037;
    value[6130] = 17'd48022;
    value[6131] = 17'd48007;
    value[6132] = 17'd47991;
    value[6133] = 17'd47976;
    value[6134] = 17'd47961;
    value[6135] = 17'd47945;
    value[6136] = 17'd47930;
    value[6137] = 17'd47915;
    value[6138] = 17'd47899;
    value[6139] = 17'd47884;
    value[6140] = 17'd47869;
    value[6141] = 17'd47853;
    value[6142] = 17'd47838;
    value[6143] = 17'd47823;
    value[6144] = 17'd47807;
    value[6145] = 17'd47792;
    value[6146] = 17'd47777;
    value[6147] = 17'd47761;
    value[6148] = 17'd47746;
    value[6149] = 17'd47731;
    value[6150] = 17'd47715;
    value[6151] = 17'd47700;
    value[6152] = 17'd47685;
    value[6153] = 17'd47669;
    value[6154] = 17'd47654;
    value[6155] = 17'd47639;
    value[6156] = 17'd47623;
    value[6157] = 17'd47608;
    value[6158] = 17'd47593;
    value[6159] = 17'd47577;
    value[6160] = 17'd47562;
    value[6161] = 17'd47547;
    value[6162] = 17'd47531;
    value[6163] = 17'd47516;
    value[6164] = 17'd47501;
    value[6165] = 17'd47485;
    value[6166] = 17'd47470;
    value[6167] = 17'd47454;
    value[6168] = 17'd47439;
    value[6169] = 17'd47424;
    value[6170] = 17'd47408;
    value[6171] = 17'd47393;
    value[6172] = 17'd47378;
    value[6173] = 17'd47362;
    value[6174] = 17'd47347;
    value[6175] = 17'd47331;
    value[6176] = 17'd47316;
    value[6177] = 17'd47301;
    value[6178] = 17'd47285;
    value[6179] = 17'd47270;
    value[6180] = 17'd47255;
    value[6181] = 17'd47239;
    value[6182] = 17'd47224;
    value[6183] = 17'd47208;
    value[6184] = 17'd47193;
    value[6185] = 17'd47178;
    value[6186] = 17'd47162;
    value[6187] = 17'd47147;
    value[6188] = 17'd47131;
    value[6189] = 17'd47116;
    value[6190] = 17'd47101;
    value[6191] = 17'd47085;
    value[6192] = 17'd47070;
    value[6193] = 17'd47054;
    value[6194] = 17'd47039;
    value[6195] = 17'd47024;
    value[6196] = 17'd47008;
    value[6197] = 17'd46993;
    value[6198] = 17'd46977;
    value[6199] = 17'd46962;
    value[6200] = 17'd46947;
    value[6201] = 17'd46931;
    value[6202] = 17'd46916;
    value[6203] = 17'd46900;
    value[6204] = 17'd46885;
    value[6205] = 17'd46870;
    value[6206] = 17'd46854;
    value[6207] = 17'd46839;
    value[6208] = 17'd46823;
    value[6209] = 17'd46808;
    value[6210] = 17'd46792;
    value[6211] = 17'd46777;
    value[6212] = 17'd46762;
    value[6213] = 17'd46746;
    value[6214] = 17'd46731;
    value[6215] = 17'd46715;
    value[6216] = 17'd46700;
    value[6217] = 17'd46684;
    value[6218] = 17'd46669;
    value[6219] = 17'd46654;
    value[6220] = 17'd46638;
    value[6221] = 17'd46623;
    value[6222] = 17'd46607;
    value[6223] = 17'd46592;
    value[6224] = 17'd46576;
    value[6225] = 17'd46561;
    value[6226] = 17'd46546;
    value[6227] = 17'd46530;
    value[6228] = 17'd46515;
    value[6229] = 17'd46499;
    value[6230] = 17'd46484;
    value[6231] = 17'd46468;
    value[6232] = 17'd46453;
    value[6233] = 17'd46437;
    value[6234] = 17'd46422;
    value[6235] = 17'd46406;
    value[6236] = 17'd46391;
    value[6237] = 17'd46376;
    value[6238] = 17'd46360;
    value[6239] = 17'd46345;
    value[6240] = 17'd46329;
    value[6241] = 17'd46314;
    value[6242] = 17'd46298;
    value[6243] = 17'd46283;
    value[6244] = 17'd46267;
    value[6245] = 17'd46252;
    value[6246] = 17'd46236;
    value[6247] = 17'd46221;
    value[6248] = 17'd46205;
    value[6249] = 17'd46190;
    value[6250] = 17'd46174;
    value[6251] = 17'd46159;
    value[6252] = 17'd46143;
    value[6253] = 17'd46128;
    value[6254] = 17'd46112;
    value[6255] = 17'd46097;
    value[6256] = 17'd46081;
    value[6257] = 17'd46066;
    value[6258] = 17'd46050;
    value[6259] = 17'd46035;
    value[6260] = 17'd46019;
    value[6261] = 17'd46004;
    value[6262] = 17'd45988;
    value[6263] = 17'd45973;
    value[6264] = 17'd45957;
    value[6265] = 17'd45942;
    value[6266] = 17'd45926;
    value[6267] = 17'd45911;
    value[6268] = 17'd45895;
    value[6269] = 17'd45880;
    value[6270] = 17'd45864;
    value[6271] = 17'd45849;
    value[6272] = 17'd45833;
    value[6273] = 17'd45818;
    value[6274] = 17'd45802;
    value[6275] = 17'd45787;
    value[6276] = 17'd45771;
    value[6277] = 17'd45756;
    value[6278] = 17'd45740;
    value[6279] = 17'd45725;
    value[6280] = 17'd45709;
    value[6281] = 17'd45694;
    value[6282] = 17'd45678;
    value[6283] = 17'd45663;
    value[6284] = 17'd45647;
    value[6285] = 17'd45632;
    value[6286] = 17'd45616;
    value[6287] = 17'd45601;
    value[6288] = 17'd45585;
    value[6289] = 17'd45570;
    value[6290] = 17'd45554;
    value[6291] = 17'd45538;
    value[6292] = 17'd45523;
    value[6293] = 17'd45507;
    value[6294] = 17'd45492;
    value[6295] = 17'd45476;
    value[6296] = 17'd45461;
    value[6297] = 17'd45445;
    value[6298] = 17'd45430;
    value[6299] = 17'd45414;
    value[6300] = 17'd45399;
    value[6301] = 17'd45383;
    value[6302] = 17'd45367;
    value[6303] = 17'd45352;
    value[6304] = 17'd45336;
    value[6305] = 17'd45321;
    value[6306] = 17'd45305;
    value[6307] = 17'd45290;
    value[6308] = 17'd45274;
    value[6309] = 17'd45259;
    value[6310] = 17'd45243;
    value[6311] = 17'd45227;
    value[6312] = 17'd45212;
    value[6313] = 17'd45196;
    value[6314] = 17'd45181;
    value[6315] = 17'd45165;
    value[6316] = 17'd45150;
    value[6317] = 17'd45134;
    value[6318] = 17'd45118;
    value[6319] = 17'd45103;
    value[6320] = 17'd45087;
    value[6321] = 17'd45072;
    value[6322] = 17'd45056;
    value[6323] = 17'd45041;
    value[6324] = 17'd45025;
    value[6325] = 17'd45009;
    value[6326] = 17'd44994;
    value[6327] = 17'd44978;
    value[6328] = 17'd44963;
    value[6329] = 17'd44947;
    value[6330] = 17'd44931;
    value[6331] = 17'd44916;
    value[6332] = 17'd44900;
    value[6333] = 17'd44885;
    value[6334] = 17'd44869;
    value[6335] = 17'd44853;
    value[6336] = 17'd44838;
    value[6337] = 17'd44822;
    value[6338] = 17'd44807;
    value[6339] = 17'd44791;
    value[6340] = 17'd44775;
    value[6341] = 17'd44760;
    value[6342] = 17'd44744;
    value[6343] = 17'd44729;
    value[6344] = 17'd44713;
    value[6345] = 17'd44697;
    value[6346] = 17'd44682;
    value[6347] = 17'd44666;
    value[6348] = 17'd44651;
    value[6349] = 17'd44635;
    value[6350] = 17'd44619;
    value[6351] = 17'd44604;
    value[6352] = 17'd44588;
    value[6353] = 17'd44572;
    value[6354] = 17'd44557;
    value[6355] = 17'd44541;
    value[6356] = 17'd44526;
    value[6357] = 17'd44510;
    value[6358] = 17'd44494;
    value[6359] = 17'd44479;
    value[6360] = 17'd44463;
    value[6361] = 17'd44447;
    value[6362] = 17'd44432;
    value[6363] = 17'd44416;
    value[6364] = 17'd44400;
    value[6365] = 17'd44385;
    value[6366] = 17'd44369;
    value[6367] = 17'd44354;
    value[6368] = 17'd44338;
    value[6369] = 17'd44322;
    value[6370] = 17'd44307;
    value[6371] = 17'd44291;
    value[6372] = 17'd44275;
    value[6373] = 17'd44260;
    value[6374] = 17'd44244;
    value[6375] = 17'd44228;
    value[6376] = 17'd44213;
    value[6377] = 17'd44197;
    value[6378] = 17'd44181;
    value[6379] = 17'd44166;
    value[6380] = 17'd44150;
    value[6381] = 17'd44134;
    value[6382] = 17'd44119;
    value[6383] = 17'd44103;
    value[6384] = 17'd44087;
    value[6385] = 17'd44072;
    value[6386] = 17'd44056;
    value[6387] = 17'd44040;
    value[6388] = 17'd44025;
    value[6389] = 17'd44009;
    value[6390] = 17'd43993;
    value[6391] = 17'd43978;
    value[6392] = 17'd43962;
    value[6393] = 17'd43946;
    value[6394] = 17'd43931;
    value[6395] = 17'd43915;
    value[6396] = 17'd43899;
    value[6397] = 17'd43884;
    value[6398] = 17'd43868;
    value[6399] = 17'd43852;
    value[6400] = 17'd43837;
    value[6401] = 17'd43821;
    value[6402] = 17'd43805;
    value[6403] = 17'd43790;
    value[6404] = 17'd43774;
    value[6405] = 17'd43758;
    value[6406] = 17'd43742;
    value[6407] = 17'd43727;
    value[6408] = 17'd43711;
    value[6409] = 17'd43695;
    value[6410] = 17'd43680;
    value[6411] = 17'd43664;
    value[6412] = 17'd43648;
    value[6413] = 17'd43633;
    value[6414] = 17'd43617;
    value[6415] = 17'd43601;
    value[6416] = 17'd43585;
    value[6417] = 17'd43570;
    value[6418] = 17'd43554;
    value[6419] = 17'd43538;
    value[6420] = 17'd43523;
    value[6421] = 17'd43507;
    value[6422] = 17'd43491;
    value[6423] = 17'd43475;
    value[6424] = 17'd43460;
    value[6425] = 17'd43444;
    value[6426] = 17'd43428;
    value[6427] = 17'd43413;
    value[6428] = 17'd43397;
    value[6429] = 17'd43381;
    value[6430] = 17'd43365;
    value[6431] = 17'd43350;
    value[6432] = 17'd43334;
    value[6433] = 17'd43318;
    value[6434] = 17'd43302;
    value[6435] = 17'd43287;
    value[6436] = 17'd43271;
    value[6437] = 17'd43255;
    value[6438] = 17'd43240;
    value[6439] = 17'd43224;
    value[6440] = 17'd43208;
    value[6441] = 17'd43192;
    value[6442] = 17'd43177;
    value[6443] = 17'd43161;
    value[6444] = 17'd43145;
    value[6445] = 17'd43129;
    value[6446] = 17'd43114;
    value[6447] = 17'd43098;
    value[6448] = 17'd43082;
    value[6449] = 17'd43066;
    value[6450] = 17'd43051;
    value[6451] = 17'd43035;
    value[6452] = 17'd43019;
    value[6453] = 17'd43003;
    value[6454] = 17'd42988;
    value[6455] = 17'd42972;
    value[6456] = 17'd42956;
    value[6457] = 17'd42940;
    value[6458] = 17'd42925;
    value[6459] = 17'd42909;
    value[6460] = 17'd42893;
    value[6461] = 17'd42877;
    value[6462] = 17'd42861;
    value[6463] = 17'd42846;
    value[6464] = 17'd42830;
    value[6465] = 17'd42814;
    value[6466] = 17'd42798;
    value[6467] = 17'd42783;
    value[6468] = 17'd42767;
    value[6469] = 17'd42751;
    value[6470] = 17'd42735;
    value[6471] = 17'd42720;
    value[6472] = 17'd42704;
    value[6473] = 17'd42688;
    value[6474] = 17'd42672;
    value[6475] = 17'd42656;
    value[6476] = 17'd42641;
    value[6477] = 17'd42625;
    value[6478] = 17'd42609;
    value[6479] = 17'd42593;
    value[6480] = 17'd42577;
    value[6481] = 17'd42562;
    value[6482] = 17'd42546;
    value[6483] = 17'd42530;
    value[6484] = 17'd42514;
    value[6485] = 17'd42498;
    value[6486] = 17'd42483;
    value[6487] = 17'd42467;
    value[6488] = 17'd42451;
    value[6489] = 17'd42435;
    value[6490] = 17'd42419;
    value[6491] = 17'd42404;
    value[6492] = 17'd42388;
    value[6493] = 17'd42372;
    value[6494] = 17'd42356;
    value[6495] = 17'd42340;
    value[6496] = 17'd42325;
    value[6497] = 17'd42309;
    value[6498] = 17'd42293;
    value[6499] = 17'd42277;
    value[6500] = 17'd42261;
    value[6501] = 17'd42246;
    value[6502] = 17'd42230;
    value[6503] = 17'd42214;
    value[6504] = 17'd42198;
    value[6505] = 17'd42182;
    value[6506] = 17'd42166;
    value[6507] = 17'd42151;
    value[6508] = 17'd42135;
    value[6509] = 17'd42119;
    value[6510] = 17'd42103;
    value[6511] = 17'd42087;
    value[6512] = 17'd42071;
    value[6513] = 17'd42056;
    value[6514] = 17'd42040;
    value[6515] = 17'd42024;
    value[6516] = 17'd42008;
    value[6517] = 17'd41992;
    value[6518] = 17'd41976;
    value[6519] = 17'd41961;
    value[6520] = 17'd41945;
    value[6521] = 17'd41929;
    value[6522] = 17'd41913;
    value[6523] = 17'd41897;
    value[6524] = 17'd41881;
    value[6525] = 17'd41865;
    value[6526] = 17'd41850;
    value[6527] = 17'd41834;
    value[6528] = 17'd41818;
    value[6529] = 17'd41802;
    value[6530] = 17'd41786;
    value[6531] = 17'd41770;
    value[6532] = 17'd41754;
    value[6533] = 17'd41739;
    value[6534] = 17'd41723;
    value[6535] = 17'd41707;
    value[6536] = 17'd41691;
    value[6537] = 17'd41675;
    value[6538] = 17'd41659;
    value[6539] = 17'd41643;
    value[6540] = 17'd41628;
    value[6541] = 17'd41612;
    value[6542] = 17'd41596;
    value[6543] = 17'd41580;
    value[6544] = 17'd41564;
    value[6545] = 17'd41548;
    value[6546] = 17'd41532;
    value[6547] = 17'd41516;
    value[6548] = 17'd41501;
    value[6549] = 17'd41485;
    value[6550] = 17'd41469;
    value[6551] = 17'd41453;
    value[6552] = 17'd41437;
    value[6553] = 17'd41421;
    value[6554] = 17'd41405;
    value[6555] = 17'd41389;
    value[6556] = 17'd41374;
    value[6557] = 17'd41358;
    value[6558] = 17'd41342;
    value[6559] = 17'd41326;
    value[6560] = 17'd41310;
    value[6561] = 17'd41294;
    value[6562] = 17'd41278;
    value[6563] = 17'd41262;
    value[6564] = 17'd41246;
    value[6565] = 17'd41230;
    value[6566] = 17'd41215;
    value[6567] = 17'd41199;
    value[6568] = 17'd41183;
    value[6569] = 17'd41167;
    value[6570] = 17'd41151;
    value[6571] = 17'd41135;
    value[6572] = 17'd41119;
    value[6573] = 17'd41103;
    value[6574] = 17'd41087;
    value[6575] = 17'd41071;
    value[6576] = 17'd41055;
    value[6577] = 17'd41040;
    value[6578] = 17'd41024;
    value[6579] = 17'd41008;
    value[6580] = 17'd40992;
    value[6581] = 17'd40976;
    value[6582] = 17'd40960;
    value[6583] = 17'd40944;
    value[6584] = 17'd40928;
    value[6585] = 17'd40912;
    value[6586] = 17'd40896;
    value[6587] = 17'd40880;
    value[6588] = 17'd40864;
    value[6589] = 17'd40848;
    value[6590] = 17'd40833;
    value[6591] = 17'd40817;
    value[6592] = 17'd40801;
    value[6593] = 17'd40785;
    value[6594] = 17'd40769;
    value[6595] = 17'd40753;
    value[6596] = 17'd40737;
    value[6597] = 17'd40721;
    value[6598] = 17'd40705;
    value[6599] = 17'd40689;
    value[6600] = 17'd40673;
    value[6601] = 17'd40657;
    value[6602] = 17'd40641;
    value[6603] = 17'd40625;
    value[6604] = 17'd40609;
    value[6605] = 17'd40593;
    value[6606] = 17'd40577;
    value[6607] = 17'd40562;
    value[6608] = 17'd40546;
    value[6609] = 17'd40530;
    value[6610] = 17'd40514;
    value[6611] = 17'd40498;
    value[6612] = 17'd40482;
    value[6613] = 17'd40466;
    value[6614] = 17'd40450;
    value[6615] = 17'd40434;
    value[6616] = 17'd40418;
    value[6617] = 17'd40402;
    value[6618] = 17'd40386;
    value[6619] = 17'd40370;
    value[6620] = 17'd40354;
    value[6621] = 17'd40338;
    value[6622] = 17'd40322;
    value[6623] = 17'd40306;
    value[6624] = 17'd40290;
    value[6625] = 17'd40274;
    value[6626] = 17'd40258;
    value[6627] = 17'd40242;
    value[6628] = 17'd40226;
    value[6629] = 17'd40210;
    value[6630] = 17'd40194;
    value[6631] = 17'd40178;
    value[6632] = 17'd40162;
    value[6633] = 17'd40146;
    value[6634] = 17'd40130;
    value[6635] = 17'd40114;
    value[6636] = 17'd40098;
    value[6637] = 17'd40082;
    value[6638] = 17'd40066;
    value[6639] = 17'd40050;
    value[6640] = 17'd40034;
    value[6641] = 17'd40018;
    value[6642] = 17'd40002;
    value[6643] = 17'd39986;
    value[6644] = 17'd39970;
    value[6645] = 17'd39954;
    value[6646] = 17'd39938;
    value[6647] = 17'd39922;
    value[6648] = 17'd39906;
    value[6649] = 17'd39890;
    value[6650] = 17'd39874;
    value[6651] = 17'd39858;
    value[6652] = 17'd39842;
    value[6653] = 17'd39826;
    value[6654] = 17'd39810;
    value[6655] = 17'd39794;
    value[6656] = 17'd39778;
    value[6657] = 17'd39762;
    value[6658] = 17'd39746;
    value[6659] = 17'd39730;
    value[6660] = 17'd39714;
    value[6661] = 17'd39698;
    value[6662] = 17'd39682;
    value[6663] = 17'd39666;
    value[6664] = 17'd39650;
    value[6665] = 17'd39634;
    value[6666] = 17'd39618;
    value[6667] = 17'd39602;
    value[6668] = 17'd39586;
    value[6669] = 17'd39570;
    value[6670] = 17'd39554;
    value[6671] = 17'd39538;
    value[6672] = 17'd39522;
    value[6673] = 17'd39506;
    value[6674] = 17'd39490;
    value[6675] = 17'd39474;
    value[6676] = 17'd39458;
    value[6677] = 17'd39442;
    value[6678] = 17'd39426;
    value[6679] = 17'd39410;
    value[6680] = 17'd39394;
    value[6681] = 17'd39378;
    value[6682] = 17'd39362;
    value[6683] = 17'd39346;
    value[6684] = 17'd39330;
    value[6685] = 17'd39313;
    value[6686] = 17'd39297;
    value[6687] = 17'd39281;
    value[6688] = 17'd39265;
    value[6689] = 17'd39249;
    value[6690] = 17'd39233;
    value[6691] = 17'd39217;
    value[6692] = 17'd39201;
    value[6693] = 17'd39185;
    value[6694] = 17'd39169;
    value[6695] = 17'd39153;
    value[6696] = 17'd39137;
    value[6697] = 17'd39121;
    value[6698] = 17'd39105;
    value[6699] = 17'd39089;
    value[6700] = 17'd39073;
    value[6701] = 17'd39057;
    value[6702] = 17'd39040;
    value[6703] = 17'd39024;
    value[6704] = 17'd39008;
    value[6705] = 17'd38992;
    value[6706] = 17'd38976;
    value[6707] = 17'd38960;
    value[6708] = 17'd38944;
    value[6709] = 17'd38928;
    value[6710] = 17'd38912;
    value[6711] = 17'd38896;
    value[6712] = 17'd38880;
    value[6713] = 17'd38864;
    value[6714] = 17'd38848;
    value[6715] = 17'd38831;
    value[6716] = 17'd38815;
    value[6717] = 17'd38799;
    value[6718] = 17'd38783;
    value[6719] = 17'd38767;
    value[6720] = 17'd38751;
    value[6721] = 17'd38735;
    value[6722] = 17'd38719;
    value[6723] = 17'd38703;
    value[6724] = 17'd38687;
    value[6725] = 17'd38671;
    value[6726] = 17'd38655;
    value[6727] = 17'd38638;
    value[6728] = 17'd38622;
    value[6729] = 17'd38606;
    value[6730] = 17'd38590;
    value[6731] = 17'd38574;
    value[6732] = 17'd38558;
    value[6733] = 17'd38542;
    value[6734] = 17'd38526;
    value[6735] = 17'd38510;
    value[6736] = 17'd38493;
    value[6737] = 17'd38477;
    value[6738] = 17'd38461;
    value[6739] = 17'd38445;
    value[6740] = 17'd38429;
    value[6741] = 17'd38413;
    value[6742] = 17'd38397;
    value[6743] = 17'd38381;
    value[6744] = 17'd38365;
    value[6745] = 17'd38348;
    value[6746] = 17'd38332;
    value[6747] = 17'd38316;
    value[6748] = 17'd38300;
    value[6749] = 17'd38284;
    value[6750] = 17'd38268;
    value[6751] = 17'd38252;
    value[6752] = 17'd38236;
    value[6753] = 17'd38219;
    value[6754] = 17'd38203;
    value[6755] = 17'd38187;
    value[6756] = 17'd38171;
    value[6757] = 17'd38155;
    value[6758] = 17'd38139;
    value[6759] = 17'd38123;
    value[6760] = 17'd38107;
    value[6761] = 17'd38090;
    value[6762] = 17'd38074;
    value[6763] = 17'd38058;
    value[6764] = 17'd38042;
    value[6765] = 17'd38026;
    value[6766] = 17'd38010;
    value[6767] = 17'd37994;
    value[6768] = 17'd37977;
    value[6769] = 17'd37961;
    value[6770] = 17'd37945;
    value[6771] = 17'd37929;
    value[6772] = 17'd37913;
    value[6773] = 17'd37897;
    value[6774] = 17'd37881;
    value[6775] = 17'd37864;
    value[6776] = 17'd37848;
    value[6777] = 17'd37832;
    value[6778] = 17'd37816;
    value[6779] = 17'd37800;
    value[6780] = 17'd37784;
    value[6781] = 17'd37767;
    value[6782] = 17'd37751;
    value[6783] = 17'd37735;
    value[6784] = 17'd37719;
    value[6785] = 17'd37703;
    value[6786] = 17'd37687;
    value[6787] = 17'd37670;
    value[6788] = 17'd37654;
    value[6789] = 17'd37638;
    value[6790] = 17'd37622;
    value[6791] = 17'd37606;
    value[6792] = 17'd37590;
    value[6793] = 17'd37573;
    value[6794] = 17'd37557;
    value[6795] = 17'd37541;
    value[6796] = 17'd37525;
    value[6797] = 17'd37509;
    value[6798] = 17'd37493;
    value[6799] = 17'd37476;
    value[6800] = 17'd37460;
    value[6801] = 17'd37444;
    value[6802] = 17'd37428;
    value[6803] = 17'd37412;
    value[6804] = 17'd37395;
    value[6805] = 17'd37379;
    value[6806] = 17'd37363;
    value[6807] = 17'd37347;
    value[6808] = 17'd37331;
    value[6809] = 17'd37314;
    value[6810] = 17'd37298;
    value[6811] = 17'd37282;
    value[6812] = 17'd37266;
    value[6813] = 17'd37250;
    value[6814] = 17'd37233;
    value[6815] = 17'd37217;
    value[6816] = 17'd37201;
    value[6817] = 17'd37185;
    value[6818] = 17'd37169;
    value[6819] = 17'd37152;
    value[6820] = 17'd37136;
    value[6821] = 17'd37120;
    value[6822] = 17'd37104;
    value[6823] = 17'd37088;
    value[6824] = 17'd37071;
    value[6825] = 17'd37055;
    value[6826] = 17'd37039;
    value[6827] = 17'd37023;
    value[6828] = 17'd37007;
    value[6829] = 17'd36990;
    value[6830] = 17'd36974;
    value[6831] = 17'd36958;
    value[6832] = 17'd36942;
    value[6833] = 17'd36926;
    value[6834] = 17'd36909;
    value[6835] = 17'd36893;
    value[6836] = 17'd36877;
    value[6837] = 17'd36861;
    value[6838] = 17'd36844;
    value[6839] = 17'd36828;
    value[6840] = 17'd36812;
    value[6841] = 17'd36796;
    value[6842] = 17'd36779;
    value[6843] = 17'd36763;
    value[6844] = 17'd36747;
    value[6845] = 17'd36731;
    value[6846] = 17'd36715;
    value[6847] = 17'd36698;
    value[6848] = 17'd36682;
    value[6849] = 17'd36666;
    value[6850] = 17'd36650;
    value[6851] = 17'd36633;
    value[6852] = 17'd36617;
    value[6853] = 17'd36601;
    value[6854] = 17'd36585;
    value[6855] = 17'd36568;
    value[6856] = 17'd36552;
    value[6857] = 17'd36536;
    value[6858] = 17'd36520;
    value[6859] = 17'd36503;
    value[6860] = 17'd36487;
    value[6861] = 17'd36471;
    value[6862] = 17'd36455;
    value[6863] = 17'd36438;
    value[6864] = 17'd36422;
    value[6865] = 17'd36406;
    value[6866] = 17'd36390;
    value[6867] = 17'd36373;
    value[6868] = 17'd36357;
    value[6869] = 17'd36341;
    value[6870] = 17'd36325;
    value[6871] = 17'd36308;
    value[6872] = 17'd36292;
    value[6873] = 17'd36276;
    value[6874] = 17'd36260;
    value[6875] = 17'd36243;
    value[6876] = 17'd36227;
    value[6877] = 17'd36211;
    value[6878] = 17'd36195;
    value[6879] = 17'd36178;
    value[6880] = 17'd36162;
    value[6881] = 17'd36146;
    value[6882] = 17'd36129;
    value[6883] = 17'd36113;
    value[6884] = 17'd36097;
    value[6885] = 17'd36081;
    value[6886] = 17'd36064;
    value[6887] = 17'd36048;
    value[6888] = 17'd36032;
    value[6889] = 17'd36015;
    value[6890] = 17'd35999;
    value[6891] = 17'd35983;
    value[6892] = 17'd35967;
    value[6893] = 17'd35950;
    value[6894] = 17'd35934;
    value[6895] = 17'd35918;
    value[6896] = 17'd35901;
    value[6897] = 17'd35885;
    value[6898] = 17'd35869;
    value[6899] = 17'd35853;
    value[6900] = 17'd35836;
    value[6901] = 17'd35820;
    value[6902] = 17'd35804;
    value[6903] = 17'd35787;
    value[6904] = 17'd35771;
    value[6905] = 17'd35755;
    value[6906] = 17'd35739;
    value[6907] = 17'd35722;
    value[6908] = 17'd35706;
    value[6909] = 17'd35690;
    value[6910] = 17'd35673;
    value[6911] = 17'd35657;
    value[6912] = 17'd35641;
    value[6913] = 17'd35624;
    value[6914] = 17'd35608;
    value[6915] = 17'd35592;
    value[6916] = 17'd35575;
    value[6917] = 17'd35559;
    value[6918] = 17'd35543;
    value[6919] = 17'd35527;
    value[6920] = 17'd35510;
    value[6921] = 17'd35494;
    value[6922] = 17'd35478;
    value[6923] = 17'd35461;
    value[6924] = 17'd35445;
    value[6925] = 17'd35429;
    value[6926] = 17'd35412;
    value[6927] = 17'd35396;
    value[6928] = 17'd35380;
    value[6929] = 17'd35363;
    value[6930] = 17'd35347;
    value[6931] = 17'd35331;
    value[6932] = 17'd35314;
    value[6933] = 17'd35298;
    value[6934] = 17'd35282;
    value[6935] = 17'd35265;
    value[6936] = 17'd35249;
    value[6937] = 17'd35233;
    value[6938] = 17'd35216;
    value[6939] = 17'd35200;
    value[6940] = 17'd35184;
    value[6941] = 17'd35167;
    value[6942] = 17'd35151;
    value[6943] = 17'd35135;
    value[6944] = 17'd35118;
    value[6945] = 17'd35102;
    value[6946] = 17'd35086;
    value[6947] = 17'd35069;
    value[6948] = 17'd35053;
    value[6949] = 17'd35037;
    value[6950] = 17'd35020;
    value[6951] = 17'd35004;
    value[6952] = 17'd34988;
    value[6953] = 17'd34971;
    value[6954] = 17'd34955;
    value[6955] = 17'd34938;
    value[6956] = 17'd34922;
    value[6957] = 17'd34906;
    value[6958] = 17'd34889;
    value[6959] = 17'd34873;
    value[6960] = 17'd34857;
    value[6961] = 17'd34840;
    value[6962] = 17'd34824;
    value[6963] = 17'd34808;
    value[6964] = 17'd34791;
    value[6965] = 17'd34775;
    value[6966] = 17'd34759;
    value[6967] = 17'd34742;
    value[6968] = 17'd34726;
    value[6969] = 17'd34709;
    value[6970] = 17'd34693;
    value[6971] = 17'd34677;
    value[6972] = 17'd34660;
    value[6973] = 17'd34644;
    value[6974] = 17'd34628;
    value[6975] = 17'd34611;
    value[6976] = 17'd34595;
    value[6977] = 17'd34578;
    value[6978] = 17'd34562;
    value[6979] = 17'd34546;
    value[6980] = 17'd34529;
    value[6981] = 17'd34513;
    value[6982] = 17'd34497;
    value[6983] = 17'd34480;
    value[6984] = 17'd34464;
    value[6985] = 17'd34447;
    value[6986] = 17'd34431;
    value[6987] = 17'd34415;
    value[6988] = 17'd34398;
    value[6989] = 17'd34382;
    value[6990] = 17'd34365;
    value[6991] = 17'd34349;
    value[6992] = 17'd34333;
    value[6993] = 17'd34316;
    value[6994] = 17'd34300;
    value[6995] = 17'd34284;
    value[6996] = 17'd34267;
    value[6997] = 17'd34251;
    value[6998] = 17'd34234;
    value[6999] = 17'd34218;
    value[7000] = 17'd34202;
    value[7001] = 17'd34185;
    value[7002] = 17'd34169;
    value[7003] = 17'd34152;
    value[7004] = 17'd34136;
    value[7005] = 17'd34119;
    value[7006] = 17'd34103;
    value[7007] = 17'd34087;
    value[7008] = 17'd34070;
    value[7009] = 17'd34054;
    value[7010] = 17'd34037;
    value[7011] = 17'd34021;
    value[7012] = 17'd34005;
    value[7013] = 17'd33988;
    value[7014] = 17'd33972;
    value[7015] = 17'd33955;
    value[7016] = 17'd33939;
    value[7017] = 17'd33923;
    value[7018] = 17'd33906;
    value[7019] = 17'd33890;
    value[7020] = 17'd33873;
    value[7021] = 17'd33857;
    value[7022] = 17'd33840;
    value[7023] = 17'd33824;
    value[7024] = 17'd33808;
    value[7025] = 17'd33791;
    value[7026] = 17'd33775;
    value[7027] = 17'd33758;
    value[7028] = 17'd33742;
    value[7029] = 17'd33725;
    value[7030] = 17'd33709;
    value[7031] = 17'd33693;
    value[7032] = 17'd33676;
    value[7033] = 17'd33660;
    value[7034] = 17'd33643;
    value[7035] = 17'd33627;
    value[7036] = 17'd33610;
    value[7037] = 17'd33594;
    value[7038] = 17'd33578;
    value[7039] = 17'd33561;
    value[7040] = 17'd33545;
    value[7041] = 17'd33528;
    value[7042] = 17'd33512;
    value[7043] = 17'd33495;
    value[7044] = 17'd33479;
    value[7045] = 17'd33462;
    value[7046] = 17'd33446;
    value[7047] = 17'd33430;
    value[7048] = 17'd33413;
    value[7049] = 17'd33397;
    value[7050] = 17'd33380;
    value[7051] = 17'd33364;
    value[7052] = 17'd33347;
    value[7053] = 17'd33331;
    value[7054] = 17'd33314;
    value[7055] = 17'd33298;
    value[7056] = 17'd33281;
    value[7057] = 17'd33265;
    value[7058] = 17'd33249;
    value[7059] = 17'd33232;
    value[7060] = 17'd33216;
    value[7061] = 17'd33199;
    value[7062] = 17'd33183;
    value[7063] = 17'd33166;
    value[7064] = 17'd33150;
    value[7065] = 17'd33133;
    value[7066] = 17'd33117;
    value[7067] = 17'd33100;
    value[7068] = 17'd33084;
    value[7069] = 17'd33067;
    value[7070] = 17'd33051;
    value[7071] = 17'd33034;
    value[7072] = 17'd33018;
    value[7073] = 17'd33002;
    value[7074] = 17'd32985;
    value[7075] = 17'd32969;
    value[7076] = 17'd32952;
    value[7077] = 17'd32936;
    value[7078] = 17'd32919;
    value[7079] = 17'd32903;
    value[7080] = 17'd32886;
    value[7081] = 17'd32870;
    value[7082] = 17'd32853;
    value[7083] = 17'd32837;
    value[7084] = 17'd32820;
    value[7085] = 17'd32804;
    value[7086] = 17'd32787;
    value[7087] = 17'd32771;
    value[7088] = 17'd32754;
    value[7089] = 17'd32738;
    value[7090] = 17'd32721;
    value[7091] = 17'd32705;
    value[7092] = 17'd32688;
    value[7093] = 17'd32672;
    value[7094] = 17'd32655;
    value[7095] = 17'd32639;
    value[7096] = 17'd32622;
    value[7097] = 17'd32606;
    value[7098] = 17'd32589;
    value[7099] = 17'd32573;
    value[7100] = 17'd32556;
    value[7101] = 17'd32540;
    value[7102] = 17'd32523;
    value[7103] = 17'd32507;
    value[7104] = 17'd32490;
    value[7105] = 17'd32474;
    value[7106] = 17'd32457;
    value[7107] = 17'd32441;
    value[7108] = 17'd32424;
    value[7109] = 17'd32408;
    value[7110] = 17'd32391;
    value[7111] = 17'd32375;
    value[7112] = 17'd32358;
    value[7113] = 17'd32342;
    value[7114] = 17'd32325;
    value[7115] = 17'd32309;
    value[7116] = 17'd32292;
    value[7117] = 17'd32276;
    value[7118] = 17'd32259;
    value[7119] = 17'd32243;
    value[7120] = 17'd32226;
    value[7121] = 17'd32210;
    value[7122] = 17'd32193;
    value[7123] = 17'd32176;
    value[7124] = 17'd32160;
    value[7125] = 17'd32143;
    value[7126] = 17'd32127;
    value[7127] = 17'd32110;
    value[7128] = 17'd32094;
    value[7129] = 17'd32077;
    value[7130] = 17'd32061;
    value[7131] = 17'd32044;
    value[7132] = 17'd32028;
    value[7133] = 17'd32011;
    value[7134] = 17'd31995;
    value[7135] = 17'd31978;
    value[7136] = 17'd31962;
    value[7137] = 17'd31945;
    value[7138] = 17'd31929;
    value[7139] = 17'd31912;
    value[7140] = 17'd31895;
    value[7141] = 17'd31879;
    value[7142] = 17'd31862;
    value[7143] = 17'd31846;
    value[7144] = 17'd31829;
    value[7145] = 17'd31813;
    value[7146] = 17'd31796;
    value[7147] = 17'd31780;
    value[7148] = 17'd31763;
    value[7149] = 17'd31747;
    value[7150] = 17'd31730;
    value[7151] = 17'd31713;
    value[7152] = 17'd31697;
    value[7153] = 17'd31680;
    value[7154] = 17'd31664;
    value[7155] = 17'd31647;
    value[7156] = 17'd31631;
    value[7157] = 17'd31614;
    value[7158] = 17'd31598;
    value[7159] = 17'd31581;
    value[7160] = 17'd31564;
    value[7161] = 17'd31548;
    value[7162] = 17'd31531;
    value[7163] = 17'd31515;
    value[7164] = 17'd31498;
    value[7165] = 17'd31482;
    value[7166] = 17'd31465;
    value[7167] = 17'd31448;
    value[7168] = 17'd31432;
    value[7169] = 17'd31415;
    value[7170] = 17'd31399;
    value[7171] = 17'd31382;
    value[7172] = 17'd31366;
    value[7173] = 17'd31349;
    value[7174] = 17'd31332;
    value[7175] = 17'd31316;
    value[7176] = 17'd31299;
    value[7177] = 17'd31283;
    value[7178] = 17'd31266;
    value[7179] = 17'd31250;
    value[7180] = 17'd31233;
    value[7181] = 17'd31216;
    value[7182] = 17'd31200;
    value[7183] = 17'd31183;
    value[7184] = 17'd31167;
    value[7185] = 17'd31150;
    value[7186] = 17'd31133;
    value[7187] = 17'd31117;
    value[7188] = 17'd31100;
    value[7189] = 17'd31084;
    value[7190] = 17'd31067;
    value[7191] = 17'd31051;
    value[7192] = 17'd31034;
    value[7193] = 17'd31017;
    value[7194] = 17'd31001;
    value[7195] = 17'd30984;
    value[7196] = 17'd30968;
    value[7197] = 17'd30951;
    value[7198] = 17'd30934;
    value[7199] = 17'd30918;
    value[7200] = 17'd30901;
    value[7201] = 17'd30885;
    value[7202] = 17'd30868;
    value[7203] = 17'd30851;
    value[7204] = 17'd30835;
    value[7205] = 17'd30818;
    value[7206] = 17'd30802;
    value[7207] = 17'd30785;
    value[7208] = 17'd30768;
    value[7209] = 17'd30752;
    value[7210] = 17'd30735;
    value[7211] = 17'd30719;
    value[7212] = 17'd30702;
    value[7213] = 17'd30685;
    value[7214] = 17'd30669;
    value[7215] = 17'd30652;
    value[7216] = 17'd30635;
    value[7217] = 17'd30619;
    value[7218] = 17'd30602;
    value[7219] = 17'd30586;
    value[7220] = 17'd30569;
    value[7221] = 17'd30552;
    value[7222] = 17'd30536;
    value[7223] = 17'd30519;
    value[7224] = 17'd30503;
    value[7225] = 17'd30486;
    value[7226] = 17'd30469;
    value[7227] = 17'd30453;
    value[7228] = 17'd30436;
    value[7229] = 17'd30419;
    value[7230] = 17'd30403;
    value[7231] = 17'd30386;
    value[7232] = 17'd30370;
    value[7233] = 17'd30353;
    value[7234] = 17'd30336;
    value[7235] = 17'd30320;
    value[7236] = 17'd30303;
    value[7237] = 17'd30286;
    value[7238] = 17'd30270;
    value[7239] = 17'd30253;
    value[7240] = 17'd30236;
    value[7241] = 17'd30220;
    value[7242] = 17'd30203;
    value[7243] = 17'd30187;
    value[7244] = 17'd30170;
    value[7245] = 17'd30153;
    value[7246] = 17'd30137;
    value[7247] = 17'd30120;
    value[7248] = 17'd30103;
    value[7249] = 17'd30087;
    value[7250] = 17'd30070;
    value[7251] = 17'd30053;
    value[7252] = 17'd30037;
    value[7253] = 17'd30020;
    value[7254] = 17'd30003;
    value[7255] = 17'd29987;
    value[7256] = 17'd29970;
    value[7257] = 17'd29954;
    value[7258] = 17'd29937;
    value[7259] = 17'd29920;
    value[7260] = 17'd29904;
    value[7261] = 17'd29887;
    value[7262] = 17'd29870;
    value[7263] = 17'd29854;
    value[7264] = 17'd29837;
    value[7265] = 17'd29820;
    value[7266] = 17'd29804;
    value[7267] = 17'd29787;
    value[7268] = 17'd29770;
    value[7269] = 17'd29754;
    value[7270] = 17'd29737;
    value[7271] = 17'd29720;
    value[7272] = 17'd29704;
    value[7273] = 17'd29687;
    value[7274] = 17'd29670;
    value[7275] = 17'd29654;
    value[7276] = 17'd29637;
    value[7277] = 17'd29620;
    value[7278] = 17'd29604;
    value[7279] = 17'd29587;
    value[7280] = 17'd29570;
    value[7281] = 17'd29554;
    value[7282] = 17'd29537;
    value[7283] = 17'd29520;
    value[7284] = 17'd29504;
    value[7285] = 17'd29487;
    value[7286] = 17'd29470;
    value[7287] = 17'd29454;
    value[7288] = 17'd29437;
    value[7289] = 17'd29420;
    value[7290] = 17'd29404;
    value[7291] = 17'd29387;
    value[7292] = 17'd29370;
    value[7293] = 17'd29353;
    value[7294] = 17'd29337;
    value[7295] = 17'd29320;
    value[7296] = 17'd29303;
    value[7297] = 17'd29287;
    value[7298] = 17'd29270;
    value[7299] = 17'd29253;
    value[7300] = 17'd29237;
    value[7301] = 17'd29220;
    value[7302] = 17'd29203;
    value[7303] = 17'd29187;
    value[7304] = 17'd29170;
    value[7305] = 17'd29153;
    value[7306] = 17'd29137;
    value[7307] = 17'd29120;
    value[7308] = 17'd29103;
    value[7309] = 17'd29086;
    value[7310] = 17'd29070;
    value[7311] = 17'd29053;
    value[7312] = 17'd29036;
    value[7313] = 17'd29020;
    value[7314] = 17'd29003;
    value[7315] = 17'd28986;
    value[7316] = 17'd28970;
    value[7317] = 17'd28953;
    value[7318] = 17'd28936;
    value[7319] = 17'd28919;
    value[7320] = 17'd28903;
    value[7321] = 17'd28886;
    value[7322] = 17'd28869;
    value[7323] = 17'd28853;
    value[7324] = 17'd28836;
    value[7325] = 17'd28819;
    value[7326] = 17'd28802;
    value[7327] = 17'd28786;
    value[7328] = 17'd28769;
    value[7329] = 17'd28752;
    value[7330] = 17'd28736;
    value[7331] = 17'd28719;
    value[7332] = 17'd28702;
    value[7333] = 17'd28685;
    value[7334] = 17'd28669;
    value[7335] = 17'd28652;
    value[7336] = 17'd28635;
    value[7337] = 17'd28619;
    value[7338] = 17'd28602;
    value[7339] = 17'd28585;
    value[7340] = 17'd28568;
    value[7341] = 17'd28552;
    value[7342] = 17'd28535;
    value[7343] = 17'd28518;
    value[7344] = 17'd28501;
    value[7345] = 17'd28485;
    value[7346] = 17'd28468;
    value[7347] = 17'd28451;
    value[7348] = 17'd28435;
    value[7349] = 17'd28418;
    value[7350] = 17'd28401;
    value[7351] = 17'd28384;
    value[7352] = 17'd28368;
    value[7353] = 17'd28351;
    value[7354] = 17'd28334;
    value[7355] = 17'd28317;
    value[7356] = 17'd28301;
    value[7357] = 17'd28284;
    value[7358] = 17'd28267;
    value[7359] = 17'd28250;
    value[7360] = 17'd28234;
    value[7361] = 17'd28217;
    value[7362] = 17'd28200;
    value[7363] = 17'd28183;
    value[7364] = 17'd28167;
    value[7365] = 17'd28150;
    value[7366] = 17'd28133;
    value[7367] = 17'd28116;
    value[7368] = 17'd28100;
    value[7369] = 17'd28083;
    value[7370] = 17'd28066;
    value[7371] = 17'd28049;
    value[7372] = 17'd28033;
    value[7373] = 17'd28016;
    value[7374] = 17'd27999;
    value[7375] = 17'd27982;
    value[7376] = 17'd27966;
    value[7377] = 17'd27949;
    value[7378] = 17'd27932;
    value[7379] = 17'd27915;
    value[7380] = 17'd27899;
    value[7381] = 17'd27882;
    value[7382] = 17'd27865;
    value[7383] = 17'd27848;
    value[7384] = 17'd27832;
    value[7385] = 17'd27815;
    value[7386] = 17'd27798;
    value[7387] = 17'd27781;
    value[7388] = 17'd27765;
    value[7389] = 17'd27748;
    value[7390] = 17'd27731;
    value[7391] = 17'd27714;
    value[7392] = 17'd27697;
    value[7393] = 17'd27681;
    value[7394] = 17'd27664;
    value[7395] = 17'd27647;
    value[7396] = 17'd27630;
    value[7397] = 17'd27614;
    value[7398] = 17'd27597;
    value[7399] = 17'd27580;
    value[7400] = 17'd27563;
    value[7401] = 17'd27546;
    value[7402] = 17'd27530;
    value[7403] = 17'd27513;
    value[7404] = 17'd27496;
    value[7405] = 17'd27479;
    value[7406] = 17'd27463;
    value[7407] = 17'd27446;
    value[7408] = 17'd27429;
    value[7409] = 17'd27412;
    value[7410] = 17'd27395;
    value[7411] = 17'd27379;
    value[7412] = 17'd27362;
    value[7413] = 17'd27345;
    value[7414] = 17'd27328;
    value[7415] = 17'd27311;
    value[7416] = 17'd27295;
    value[7417] = 17'd27278;
    value[7418] = 17'd27261;
    value[7419] = 17'd27244;
    value[7420] = 17'd27228;
    value[7421] = 17'd27211;
    value[7422] = 17'd27194;
    value[7423] = 17'd27177;
    value[7424] = 17'd27160;
    value[7425] = 17'd27144;
    value[7426] = 17'd27127;
    value[7427] = 17'd27110;
    value[7428] = 17'd27093;
    value[7429] = 17'd27076;
    value[7430] = 17'd27060;
    value[7431] = 17'd27043;
    value[7432] = 17'd27026;
    value[7433] = 17'd27009;
    value[7434] = 17'd26992;
    value[7435] = 17'd26976;
    value[7436] = 17'd26959;
    value[7437] = 17'd26942;
    value[7438] = 17'd26925;
    value[7439] = 17'd26908;
    value[7440] = 17'd26891;
    value[7441] = 17'd26875;
    value[7442] = 17'd26858;
    value[7443] = 17'd26841;
    value[7444] = 17'd26824;
    value[7445] = 17'd26807;
    value[7446] = 17'd26791;
    value[7447] = 17'd26774;
    value[7448] = 17'd26757;
    value[7449] = 17'd26740;
    value[7450] = 17'd26723;
    value[7451] = 17'd26707;
    value[7452] = 17'd26690;
    value[7453] = 17'd26673;
    value[7454] = 17'd26656;
    value[7455] = 17'd26639;
    value[7456] = 17'd26622;
    value[7457] = 17'd26606;
    value[7458] = 17'd26589;
    value[7459] = 17'd26572;
    value[7460] = 17'd26555;
    value[7461] = 17'd26538;
    value[7462] = 17'd26521;
    value[7463] = 17'd26505;
    value[7464] = 17'd26488;
    value[7465] = 17'd26471;
    value[7466] = 17'd26454;
    value[7467] = 17'd26437;
    value[7468] = 17'd26420;
    value[7469] = 17'd26404;
    value[7470] = 17'd26387;
    value[7471] = 17'd26370;
    value[7472] = 17'd26353;
    value[7473] = 17'd26336;
    value[7474] = 17'd26319;
    value[7475] = 17'd26303;
    value[7476] = 17'd26286;
    value[7477] = 17'd26269;
    value[7478] = 17'd26252;
    value[7479] = 17'd26235;
    value[7480] = 17'd26218;
    value[7481] = 17'd26202;
    value[7482] = 17'd26185;
    value[7483] = 17'd26168;
    value[7484] = 17'd26151;
    value[7485] = 17'd26134;
    value[7486] = 17'd26117;
    value[7487] = 17'd26101;
    value[7488] = 17'd26084;
    value[7489] = 17'd26067;
    value[7490] = 17'd26050;
    value[7491] = 17'd26033;
    value[7492] = 17'd26016;
    value[7493] = 17'd25999;
    value[7494] = 17'd25983;
    value[7495] = 17'd25966;
    value[7496] = 17'd25949;
    value[7497] = 17'd25932;
    value[7498] = 17'd25915;
    value[7499] = 17'd25898;
    value[7500] = 17'd25881;
    value[7501] = 17'd25865;
    value[7502] = 17'd25848;
    value[7503] = 17'd25831;
    value[7504] = 17'd25814;
    value[7505] = 17'd25797;
    value[7506] = 17'd25780;
    value[7507] = 17'd25763;
    value[7508] = 17'd25747;
    value[7509] = 17'd25730;
    value[7510] = 17'd25713;
    value[7511] = 17'd25696;
    value[7512] = 17'd25679;
    value[7513] = 17'd25662;
    value[7514] = 17'd25645;
    value[7515] = 17'd25628;
    value[7516] = 17'd25612;
    value[7517] = 17'd25595;
    value[7518] = 17'd25578;
    value[7519] = 17'd25561;
    value[7520] = 17'd25544;
    value[7521] = 17'd25527;
    value[7522] = 17'd25510;
    value[7523] = 17'd25493;
    value[7524] = 17'd25477;
    value[7525] = 17'd25460;
    value[7526] = 17'd25443;
    value[7527] = 17'd25426;
    value[7528] = 17'd25409;
    value[7529] = 17'd25392;
    value[7530] = 17'd25375;
    value[7531] = 17'd25358;
    value[7532] = 17'd25342;
    value[7533] = 17'd25325;
    value[7534] = 17'd25308;
    value[7535] = 17'd25291;
    value[7536] = 17'd25274;
    value[7537] = 17'd25257;
    value[7538] = 17'd25240;
    value[7539] = 17'd25223;
    value[7540] = 17'd25206;
    value[7541] = 17'd25190;
    value[7542] = 17'd25173;
    value[7543] = 17'd25156;
    value[7544] = 17'd25139;
    value[7545] = 17'd25122;
    value[7546] = 17'd25105;
    value[7547] = 17'd25088;
    value[7548] = 17'd25071;
    value[7549] = 17'd25054;
    value[7550] = 17'd25038;
    value[7551] = 17'd25021;
    value[7552] = 17'd25004;
    value[7553] = 17'd24987;
    value[7554] = 17'd24970;
    value[7555] = 17'd24953;
    value[7556] = 17'd24936;
    value[7557] = 17'd24919;
    value[7558] = 17'd24902;
    value[7559] = 17'd24885;
    value[7560] = 17'd24868;
    value[7561] = 17'd24852;
    value[7562] = 17'd24835;
    value[7563] = 17'd24818;
    value[7564] = 17'd24801;
    value[7565] = 17'd24784;
    value[7566] = 17'd24767;
    value[7567] = 17'd24750;
    value[7568] = 17'd24733;
    value[7569] = 17'd24716;
    value[7570] = 17'd24699;
    value[7571] = 17'd24682;
    value[7572] = 17'd24666;
    value[7573] = 17'd24649;
    value[7574] = 17'd24632;
    value[7575] = 17'd24615;
    value[7576] = 17'd24598;
    value[7577] = 17'd24581;
    value[7578] = 17'd24564;
    value[7579] = 17'd24547;
    value[7580] = 17'd24530;
    value[7581] = 17'd24513;
    value[7582] = 17'd24496;
    value[7583] = 17'd24479;
    value[7584] = 17'd24463;
    value[7585] = 17'd24446;
    value[7586] = 17'd24429;
    value[7587] = 17'd24412;
    value[7588] = 17'd24395;
    value[7589] = 17'd24378;
    value[7590] = 17'd24361;
    value[7591] = 17'd24344;
    value[7592] = 17'd24327;
    value[7593] = 17'd24310;
    value[7594] = 17'd24293;
    value[7595] = 17'd24276;
    value[7596] = 17'd24259;
    value[7597] = 17'd24242;
    value[7598] = 17'd24226;
    value[7599] = 17'd24209;
    value[7600] = 17'd24192;
    value[7601] = 17'd24175;
    value[7602] = 17'd24158;
    value[7603] = 17'd24141;
    value[7604] = 17'd24124;
    value[7605] = 17'd24107;
    value[7606] = 17'd24090;
    value[7607] = 17'd24073;
    value[7608] = 17'd24056;
    value[7609] = 17'd24039;
    value[7610] = 17'd24022;
    value[7611] = 17'd24005;
    value[7612] = 17'd23988;
    value[7613] = 17'd23971;
    value[7614] = 17'd23955;
    value[7615] = 17'd23938;
    value[7616] = 17'd23921;
    value[7617] = 17'd23904;
    value[7618] = 17'd23887;
    value[7619] = 17'd23870;
    value[7620] = 17'd23853;
    value[7621] = 17'd23836;
    value[7622] = 17'd23819;
    value[7623] = 17'd23802;
    value[7624] = 17'd23785;
    value[7625] = 17'd23768;
    value[7626] = 17'd23751;
    value[7627] = 17'd23734;
    value[7628] = 17'd23717;
    value[7629] = 17'd23700;
    value[7630] = 17'd23683;
    value[7631] = 17'd23666;
    value[7632] = 17'd23649;
    value[7633] = 17'd23632;
    value[7634] = 17'd23615;
    value[7635] = 17'd23599;
    value[7636] = 17'd23582;
    value[7637] = 17'd23565;
    value[7638] = 17'd23548;
    value[7639] = 17'd23531;
    value[7640] = 17'd23514;
    value[7641] = 17'd23497;
    value[7642] = 17'd23480;
    value[7643] = 17'd23463;
    value[7644] = 17'd23446;
    value[7645] = 17'd23429;
    value[7646] = 17'd23412;
    value[7647] = 17'd23395;
    value[7648] = 17'd23378;
    value[7649] = 17'd23361;
    value[7650] = 17'd23344;
    value[7651] = 17'd23327;
    value[7652] = 17'd23310;
    value[7653] = 17'd23293;
    value[7654] = 17'd23276;
    value[7655] = 17'd23259;
    value[7656] = 17'd23242;
    value[7657] = 17'd23225;
    value[7658] = 17'd23208;
    value[7659] = 17'd23191;
    value[7660] = 17'd23174;
    value[7661] = 17'd23157;
    value[7662] = 17'd23140;
    value[7663] = 17'd23123;
    value[7664] = 17'd23106;
    value[7665] = 17'd23089;
    value[7666] = 17'd23072;
    value[7667] = 17'd23055;
    value[7668] = 17'd23038;
    value[7669] = 17'd23021;
    value[7670] = 17'd23004;
    value[7671] = 17'd22987;
    value[7672] = 17'd22971;
    value[7673] = 17'd22954;
    value[7674] = 17'd22937;
    value[7675] = 17'd22920;
    value[7676] = 17'd22903;
    value[7677] = 17'd22886;
    value[7678] = 17'd22869;
    value[7679] = 17'd22852;
    value[7680] = 17'd22835;
    value[7681] = 17'd22818;
    value[7682] = 17'd22801;
    value[7683] = 17'd22784;
    value[7684] = 17'd22767;
    value[7685] = 17'd22750;
    value[7686] = 17'd22733;
    value[7687] = 17'd22716;
    value[7688] = 17'd22699;
    value[7689] = 17'd22682;
    value[7690] = 17'd22665;
    value[7691] = 17'd22648;
    value[7692] = 17'd22631;
    value[7693] = 17'd22614;
    value[7694] = 17'd22597;
    value[7695] = 17'd22580;
    value[7696] = 17'd22563;
    value[7697] = 17'd22546;
    value[7698] = 17'd22529;
    value[7699] = 17'd22512;
    value[7700] = 17'd22495;
    value[7701] = 17'd22478;
    value[7702] = 17'd22461;
    value[7703] = 17'd22444;
    value[7704] = 17'd22427;
    value[7705] = 17'd22410;
    value[7706] = 17'd22393;
    value[7707] = 17'd22376;
    value[7708] = 17'd22359;
    value[7709] = 17'd22342;
    value[7710] = 17'd22325;
    value[7711] = 17'd22307;
    value[7712] = 17'd22290;
    value[7713] = 17'd22273;
    value[7714] = 17'd22256;
    value[7715] = 17'd22239;
    value[7716] = 17'd22222;
    value[7717] = 17'd22205;
    value[7718] = 17'd22188;
    value[7719] = 17'd22171;
    value[7720] = 17'd22154;
    value[7721] = 17'd22137;
    value[7722] = 17'd22120;
    value[7723] = 17'd22103;
    value[7724] = 17'd22086;
    value[7725] = 17'd22069;
    value[7726] = 17'd22052;
    value[7727] = 17'd22035;
    value[7728] = 17'd22018;
    value[7729] = 17'd22001;
    value[7730] = 17'd21984;
    value[7731] = 17'd21967;
    value[7732] = 17'd21950;
    value[7733] = 17'd21933;
    value[7734] = 17'd21916;
    value[7735] = 17'd21899;
    value[7736] = 17'd21882;
    value[7737] = 17'd21865;
    value[7738] = 17'd21848;
    value[7739] = 17'd21831;
    value[7740] = 17'd21814;
    value[7741] = 17'd21797;
    value[7742] = 17'd21780;
    value[7743] = 17'd21763;
    value[7744] = 17'd21746;
    value[7745] = 17'd21729;
    value[7746] = 17'd21712;
    value[7747] = 17'd21695;
    value[7748] = 17'd21678;
    value[7749] = 17'd21661;
    value[7750] = 17'd21643;
    value[7751] = 17'd21626;
    value[7752] = 17'd21609;
    value[7753] = 17'd21592;
    value[7754] = 17'd21575;
    value[7755] = 17'd21558;
    value[7756] = 17'd21541;
    value[7757] = 17'd21524;
    value[7758] = 17'd21507;
    value[7759] = 17'd21490;
    value[7760] = 17'd21473;
    value[7761] = 17'd21456;
    value[7762] = 17'd21439;
    value[7763] = 17'd21422;
    value[7764] = 17'd21405;
    value[7765] = 17'd21388;
    value[7766] = 17'd21371;
    value[7767] = 17'd21354;
    value[7768] = 17'd21337;
    value[7769] = 17'd21320;
    value[7770] = 17'd21303;
    value[7771] = 17'd21285;
    value[7772] = 17'd21268;
    value[7773] = 17'd21251;
    value[7774] = 17'd21234;
    value[7775] = 17'd21217;
    value[7776] = 17'd21200;
    value[7777] = 17'd21183;
    value[7778] = 17'd21166;
    value[7779] = 17'd21149;
    value[7780] = 17'd21132;
    value[7781] = 17'd21115;
    value[7782] = 17'd21098;
    value[7783] = 17'd21081;
    value[7784] = 17'd21064;
    value[7785] = 17'd21047;
    value[7786] = 17'd21030;
    value[7787] = 17'd21013;
    value[7788] = 17'd20995;
    value[7789] = 17'd20978;
    value[7790] = 17'd20961;
    value[7791] = 17'd20944;
    value[7792] = 17'd20927;
    value[7793] = 17'd20910;
    value[7794] = 17'd20893;
    value[7795] = 17'd20876;
    value[7796] = 17'd20859;
    value[7797] = 17'd20842;
    value[7798] = 17'd20825;
    value[7799] = 17'd20808;
    value[7800] = 17'd20791;
    value[7801] = 17'd20774;
    value[7802] = 17'd20757;
    value[7803] = 17'd20739;
    value[7804] = 17'd20722;
    value[7805] = 17'd20705;
    value[7806] = 17'd20688;
    value[7807] = 17'd20671;
    value[7808] = 17'd20654;
    value[7809] = 17'd20637;
    value[7810] = 17'd20620;
    value[7811] = 17'd20603;
    value[7812] = 17'd20586;
    value[7813] = 17'd20569;
    value[7814] = 17'd20552;
    value[7815] = 17'd20535;
    value[7816] = 17'd20517;
    value[7817] = 17'd20500;
    value[7818] = 17'd20483;
    value[7819] = 17'd20466;
    value[7820] = 17'd20449;
    value[7821] = 17'd20432;
    value[7822] = 17'd20415;
    value[7823] = 17'd20398;
    value[7824] = 17'd20381;
    value[7825] = 17'd20364;
    value[7826] = 17'd20347;
    value[7827] = 17'd20329;
    value[7828] = 17'd20312;
    value[7829] = 17'd20295;
    value[7830] = 17'd20278;
    value[7831] = 17'd20261;
    value[7832] = 17'd20244;
    value[7833] = 17'd20227;
    value[7834] = 17'd20210;
    value[7835] = 17'd20193;
    value[7836] = 17'd20176;
    value[7837] = 17'd20159;
    value[7838] = 17'd20141;
    value[7839] = 17'd20124;
    value[7840] = 17'd20107;
    value[7841] = 17'd20090;
    value[7842] = 17'd20073;
    value[7843] = 17'd20056;
    value[7844] = 17'd20039;
    value[7845] = 17'd20022;
    value[7846] = 17'd20005;
    value[7847] = 17'd19988;
    value[7848] = 17'd19970;
    value[7849] = 17'd19953;
    value[7850] = 17'd19936;
    value[7851] = 17'd19919;
    value[7852] = 17'd19902;
    value[7853] = 17'd19885;
    value[7854] = 17'd19868;
    value[7855] = 17'd19851;
    value[7856] = 17'd19834;
    value[7857] = 17'd19817;
    value[7858] = 17'd19799;
    value[7859] = 17'd19782;
    value[7860] = 17'd19765;
    value[7861] = 17'd19748;
    value[7862] = 17'd19731;
    value[7863] = 17'd19714;
    value[7864] = 17'd19697;
    value[7865] = 17'd19680;
    value[7866] = 17'd19663;
    value[7867] = 17'd19645;
    value[7868] = 17'd19628;
    value[7869] = 17'd19611;
    value[7870] = 17'd19594;
    value[7871] = 17'd19577;
    value[7872] = 17'd19560;
    value[7873] = 17'd19543;
    value[7874] = 17'd19526;
    value[7875] = 17'd19509;
    value[7876] = 17'd19491;
    value[7877] = 17'd19474;
    value[7878] = 17'd19457;
    value[7879] = 17'd19440;
    value[7880] = 17'd19423;
    value[7881] = 17'd19406;
    value[7882] = 17'd19389;
    value[7883] = 17'd19372;
    value[7884] = 17'd19354;
    value[7885] = 17'd19337;
    value[7886] = 17'd19320;
    value[7887] = 17'd19303;
    value[7888] = 17'd19286;
    value[7889] = 17'd19269;
    value[7890] = 17'd19252;
    value[7891] = 17'd19235;
    value[7892] = 17'd19217;
    value[7893] = 17'd19200;
    value[7894] = 17'd19183;
    value[7895] = 17'd19166;
    value[7896] = 17'd19149;
    value[7897] = 17'd19132;
    value[7898] = 17'd19115;
    value[7899] = 17'd19098;
    value[7900] = 17'd19080;
    value[7901] = 17'd19063;
    value[7902] = 17'd19046;
    value[7903] = 17'd19029;
    value[7904] = 17'd19012;
    value[7905] = 17'd18995;
    value[7906] = 17'd18978;
    value[7907] = 17'd18960;
    value[7908] = 17'd18943;
    value[7909] = 17'd18926;
    value[7910] = 17'd18909;
    value[7911] = 17'd18892;
    value[7912] = 17'd18875;
    value[7913] = 17'd18858;
    value[7914] = 17'd18840;
    value[7915] = 17'd18823;
    value[7916] = 17'd18806;
    value[7917] = 17'd18789;
    value[7918] = 17'd18772;
    value[7919] = 17'd18755;
    value[7920] = 17'd18738;
    value[7921] = 17'd18720;
    value[7922] = 17'd18703;
    value[7923] = 17'd18686;
    value[7924] = 17'd18669;
    value[7925] = 17'd18652;
    value[7926] = 17'd18635;
    value[7927] = 17'd18618;
    value[7928] = 17'd18600;
    value[7929] = 17'd18583;
    value[7930] = 17'd18566;
    value[7931] = 17'd18549;
    value[7932] = 17'd18532;
    value[7933] = 17'd18515;
    value[7934] = 17'd18498;
    value[7935] = 17'd18480;
    value[7936] = 17'd18463;
    value[7937] = 17'd18446;
    value[7938] = 17'd18429;
    value[7939] = 17'd18412;
    value[7940] = 17'd18395;
    value[7941] = 17'd18377;
    value[7942] = 17'd18360;
    value[7943] = 17'd18343;
    value[7944] = 17'd18326;
    value[7945] = 17'd18309;
    value[7946] = 17'd18292;
    value[7947] = 17'd18275;
    value[7948] = 17'd18257;
    value[7949] = 17'd18240;
    value[7950] = 17'd18223;
    value[7951] = 17'd18206;
    value[7952] = 17'd18189;
    value[7953] = 17'd18172;
    value[7954] = 17'd18154;
    value[7955] = 17'd18137;
    value[7956] = 17'd18120;
    value[7957] = 17'd18103;
    value[7958] = 17'd18086;
    value[7959] = 17'd18069;
    value[7960] = 17'd18051;
    value[7961] = 17'd18034;
    value[7962] = 17'd18017;
    value[7963] = 17'd18000;
    value[7964] = 17'd17983;
    value[7965] = 17'd17966;
    value[7966] = 17'd17948;
    value[7967] = 17'd17931;
    value[7968] = 17'd17914;
    value[7969] = 17'd17897;
    value[7970] = 17'd17880;
    value[7971] = 17'd17863;
    value[7972] = 17'd17845;
    value[7973] = 17'd17828;
    value[7974] = 17'd17811;
    value[7975] = 17'd17794;
    value[7976] = 17'd17777;
    value[7977] = 17'd17760;
    value[7978] = 17'd17742;
    value[7979] = 17'd17725;
    value[7980] = 17'd17708;
    value[7981] = 17'd17691;
    value[7982] = 17'd17674;
    value[7983] = 17'd17656;
    value[7984] = 17'd17639;
    value[7985] = 17'd17622;
    value[7986] = 17'd17605;
    value[7987] = 17'd17588;
    value[7988] = 17'd17571;
    value[7989] = 17'd17553;
    value[7990] = 17'd17536;
    value[7991] = 17'd17519;
    value[7992] = 17'd17502;
    value[7993] = 17'd17485;
    value[7994] = 17'd17467;
    value[7995] = 17'd17450;
    value[7996] = 17'd17433;
    value[7997] = 17'd17416;
    value[7998] = 17'd17399;
    value[7999] = 17'd17382;
    value[8000] = 17'd17364;
    value[8001] = 17'd17347;
    value[8002] = 17'd17330;
    value[8003] = 17'd17313;
    value[8004] = 17'd17296;
    value[8005] = 17'd17278;
    value[8006] = 17'd17261;
    value[8007] = 17'd17244;
    value[8008] = 17'd17227;
    value[8009] = 17'd17210;
    value[8010] = 17'd17192;
    value[8011] = 17'd17175;
    value[8012] = 17'd17158;
    value[8013] = 17'd17141;
    value[8014] = 17'd17124;
    value[8015] = 17'd17106;
    value[8016] = 17'd17089;
    value[8017] = 17'd17072;
    value[8018] = 17'd17055;
    value[8019] = 17'd17038;
    value[8020] = 17'd17020;
    value[8021] = 17'd17003;
    value[8022] = 17'd16986;
    value[8023] = 17'd16969;
    value[8024] = 17'd16952;
    value[8025] = 17'd16934;
    value[8026] = 17'd16917;
    value[8027] = 17'd16900;
    value[8028] = 17'd16883;
    value[8029] = 17'd16866;
    value[8030] = 17'd16848;
    value[8031] = 17'd16831;
    value[8032] = 17'd16814;
    value[8033] = 17'd16797;
    value[8034] = 17'd16780;
    value[8035] = 17'd16762;
    value[8036] = 17'd16745;
    value[8037] = 17'd16728;
    value[8038] = 17'd16711;
    value[8039] = 17'd16694;
    value[8040] = 17'd16676;
    value[8041] = 17'd16659;
    value[8042] = 17'd16642;
    value[8043] = 17'd16625;
    value[8044] = 17'd16608;
    value[8045] = 17'd16590;
    value[8046] = 17'd16573;
    value[8047] = 17'd16556;
    value[8048] = 17'd16539;
    value[8049] = 17'd16521;
    value[8050] = 17'd16504;
    value[8051] = 17'd16487;
    value[8052] = 17'd16470;
    value[8053] = 17'd16453;
    value[8054] = 17'd16435;
    value[8055] = 17'd16418;
    value[8056] = 17'd16401;
    value[8057] = 17'd16384;
    value[8058] = 17'd16367;
    value[8059] = 17'd16349;
    value[8060] = 17'd16332;
    value[8061] = 17'd16315;
    value[8062] = 17'd16298;
    value[8063] = 17'd16280;
    value[8064] = 17'd16263;
    value[8065] = 17'd16246;
    value[8066] = 17'd16229;
    value[8067] = 17'd16212;
    value[8068] = 17'd16194;
    value[8069] = 17'd16177;
    value[8070] = 17'd16160;
    value[8071] = 17'd16143;
    value[8072] = 17'd16125;
    value[8073] = 17'd16108;
    value[8074] = 17'd16091;
    value[8075] = 17'd16074;
    value[8076] = 17'd16057;
    value[8077] = 17'd16039;
    value[8078] = 17'd16022;
    value[8079] = 17'd16005;
    value[8080] = 17'd15988;
    value[8081] = 17'd15970;
    value[8082] = 17'd15953;
    value[8083] = 17'd15936;
    value[8084] = 17'd15919;
    value[8085] = 17'd15901;
    value[8086] = 17'd15884;
    value[8087] = 17'd15867;
    value[8088] = 17'd15850;
    value[8089] = 17'd15833;
    value[8090] = 17'd15815;
    value[8091] = 17'd15798;
    value[8092] = 17'd15781;
    value[8093] = 17'd15764;
    value[8094] = 17'd15746;
    value[8095] = 17'd15729;
    value[8096] = 17'd15712;
    value[8097] = 17'd15695;
    value[8098] = 17'd15677;
    value[8099] = 17'd15660;
    value[8100] = 17'd15643;
    value[8101] = 17'd15626;
    value[8102] = 17'd15608;
    value[8103] = 17'd15591;
    value[8104] = 17'd15574;
    value[8105] = 17'd15557;
    value[8106] = 17'd15540;
    value[8107] = 17'd15522;
    value[8108] = 17'd15505;
    value[8109] = 17'd15488;
    value[8110] = 17'd15471;
    value[8111] = 17'd15453;
    value[8112] = 17'd15436;
    value[8113] = 17'd15419;
    value[8114] = 17'd15402;
    value[8115] = 17'd15384;
    value[8116] = 17'd15367;
    value[8117] = 17'd15350;
    value[8118] = 17'd15333;
    value[8119] = 17'd15315;
    value[8120] = 17'd15298;
    value[8121] = 17'd15281;
    value[8122] = 17'd15264;
    value[8123] = 17'd15246;
    value[8124] = 17'd15229;
    value[8125] = 17'd15212;
    value[8126] = 17'd15195;
    value[8127] = 17'd15177;
    value[8128] = 17'd15160;
    value[8129] = 17'd15143;
    value[8130] = 17'd15126;
    value[8131] = 17'd15108;
    value[8132] = 17'd15091;
    value[8133] = 17'd15074;
    value[8134] = 17'd15057;
    value[8135] = 17'd15039;
    value[8136] = 17'd15022;
    value[8137] = 17'd15005;
    value[8138] = 17'd14988;
    value[8139] = 17'd14970;
    value[8140] = 17'd14953;
    value[8141] = 17'd14936;
    value[8142] = 17'd14919;
    value[8143] = 17'd14901;
    value[8144] = 17'd14884;
    value[8145] = 17'd14867;
    value[8146] = 17'd14849;
    value[8147] = 17'd14832;
    value[8148] = 17'd14815;
    value[8149] = 17'd14798;
    value[8150] = 17'd14780;
    value[8151] = 17'd14763;
    value[8152] = 17'd14746;
    value[8153] = 17'd14729;
    value[8154] = 17'd14711;
    value[8155] = 17'd14694;
    value[8156] = 17'd14677;
    value[8157] = 17'd14660;
    value[8158] = 17'd14642;
    value[8159] = 17'd14625;
    value[8160] = 17'd14608;
    value[8161] = 17'd14591;
    value[8162] = 17'd14573;
    value[8163] = 17'd14556;
    value[8164] = 17'd14539;
    value[8165] = 17'd14521;
    value[8166] = 17'd14504;
    value[8167] = 17'd14487;
    value[8168] = 17'd14470;
    value[8169] = 17'd14452;
    value[8170] = 17'd14435;
    value[8171] = 17'd14418;
    value[8172] = 17'd14401;
    value[8173] = 17'd14383;
    value[8174] = 17'd14366;
    value[8175] = 17'd14349;
    value[8176] = 17'd14331;
    value[8177] = 17'd14314;
    value[8178] = 17'd14297;
    value[8179] = 17'd14280;
    value[8180] = 17'd14262;
    value[8181] = 17'd14245;
    value[8182] = 17'd14228;
    value[8183] = 17'd14211;
    value[8184] = 17'd14193;
    value[8185] = 17'd14176;
    value[8186] = 17'd14159;
    value[8187] = 17'd14141;
    value[8188] = 17'd14124;
    value[8189] = 17'd14107;
    value[8190] = 17'd14090;
    value[8191] = 17'd14072;
    value[8192] = 17'd14055;
    value[8193] = 17'd14038;
    value[8194] = 17'd14021;
    value[8195] = 17'd14003;
    value[8196] = 17'd13986;
    value[8197] = 17'd13969;
    value[8198] = 17'd13951;
    value[8199] = 17'd13934;
    value[8200] = 17'd13917;
    value[8201] = 17'd13900;
    value[8202] = 17'd13882;
    value[8203] = 17'd13865;
    value[8204] = 17'd13848;
    value[8205] = 17'd13830;
    value[8206] = 17'd13813;
    value[8207] = 17'd13796;
    value[8208] = 17'd13779;
    value[8209] = 17'd13761;
    value[8210] = 17'd13744;
    value[8211] = 17'd13727;
    value[8212] = 17'd13709;
    value[8213] = 17'd13692;
    value[8214] = 17'd13675;
    value[8215] = 17'd13658;
    value[8216] = 17'd13640;
    value[8217] = 17'd13623;
    value[8218] = 17'd13606;
    value[8219] = 17'd13588;
    value[8220] = 17'd13571;
    value[8221] = 17'd13554;
    value[8222] = 17'd13536;
    value[8223] = 17'd13519;
    value[8224] = 17'd13502;
    value[8225] = 17'd13485;
    value[8226] = 17'd13467;
    value[8227] = 17'd13450;
    value[8228] = 17'd13433;
    value[8229] = 17'd13415;
    value[8230] = 17'd13398;
    value[8231] = 17'd13381;
    value[8232] = 17'd13364;
    value[8233] = 17'd13346;
    value[8234] = 17'd13329;
    value[8235] = 17'd13312;
    value[8236] = 17'd13294;
    value[8237] = 17'd13277;
    value[8238] = 17'd13260;
    value[8239] = 17'd13242;
    value[8240] = 17'd13225;
    value[8241] = 17'd13208;
    value[8242] = 17'd13191;
    value[8243] = 17'd13173;
    value[8244] = 17'd13156;
    value[8245] = 17'd13139;
    value[8246] = 17'd13121;
    value[8247] = 17'd13104;
    value[8248] = 17'd13087;
    value[8249] = 17'd13069;
    value[8250] = 17'd13052;
    value[8251] = 17'd13035;
    value[8252] = 17'd13018;
    value[8253] = 17'd13000;
    value[8254] = 17'd12983;
    value[8255] = 17'd12966;
    value[8256] = 17'd12948;
    value[8257] = 17'd12931;
    value[8258] = 17'd12914;
    value[8259] = 17'd12896;
    value[8260] = 17'd12879;
    value[8261] = 17'd12862;
    value[8262] = 17'd12844;
    value[8263] = 17'd12827;
    value[8264] = 17'd12810;
    value[8265] = 17'd12793;
    value[8266] = 17'd12775;
    value[8267] = 17'd12758;
    value[8268] = 17'd12741;
    value[8269] = 17'd12723;
    value[8270] = 17'd12706;
    value[8271] = 17'd12689;
    value[8272] = 17'd12671;
    value[8273] = 17'd12654;
    value[8274] = 17'd12637;
    value[8275] = 17'd12619;
    value[8276] = 17'd12602;
    value[8277] = 17'd12585;
    value[8278] = 17'd12567;
    value[8279] = 17'd12550;
    value[8280] = 17'd12533;
    value[8281] = 17'd12516;
    value[8282] = 17'd12498;
    value[8283] = 17'd12481;
    value[8284] = 17'd12464;
    value[8285] = 17'd12446;
    value[8286] = 17'd12429;
    value[8287] = 17'd12412;
    value[8288] = 17'd12394;
    value[8289] = 17'd12377;
    value[8290] = 17'd12360;
    value[8291] = 17'd12342;
    value[8292] = 17'd12325;
    value[8293] = 17'd12308;
    value[8294] = 17'd12290;
    value[8295] = 17'd12273;
    value[8296] = 17'd12256;
    value[8297] = 17'd12238;
    value[8298] = 17'd12221;
    value[8299] = 17'd12204;
    value[8300] = 17'd12186;
    value[8301] = 17'd12169;
    value[8302] = 17'd12152;
    value[8303] = 17'd12134;
    value[8304] = 17'd12117;
    value[8305] = 17'd12100;
    value[8306] = 17'd12082;
    value[8307] = 17'd12065;
    value[8308] = 17'd12048;
    value[8309] = 17'd12031;
    value[8310] = 17'd12013;
    value[8311] = 17'd11996;
    value[8312] = 17'd11979;
    value[8313] = 17'd11961;
    value[8314] = 17'd11944;
    value[8315] = 17'd11927;
    value[8316] = 17'd11909;
    value[8317] = 17'd11892;
    value[8318] = 17'd11875;
    value[8319] = 17'd11857;
    value[8320] = 17'd11840;
    value[8321] = 17'd11823;
    value[8322] = 17'd11805;
    value[8323] = 17'd11788;
    value[8324] = 17'd11771;
    value[8325] = 17'd11753;
    value[8326] = 17'd11736;
    value[8327] = 17'd11719;
    value[8328] = 17'd11701;
    value[8329] = 17'd11684;
    value[8330] = 17'd11667;
    value[8331] = 17'd11649;
    value[8332] = 17'd11632;
    value[8333] = 17'd11615;
    value[8334] = 17'd11597;
    value[8335] = 17'd11580;
    value[8336] = 17'd11563;
    value[8337] = 17'd11545;
    value[8338] = 17'd11528;
    value[8339] = 17'd11511;
    value[8340] = 17'd11493;
    value[8341] = 17'd11476;
    value[8342] = 17'd11459;
    value[8343] = 17'd11441;
    value[8344] = 17'd11424;
    value[8345] = 17'd11407;
    value[8346] = 17'd11389;
    value[8347] = 17'd11372;
    value[8348] = 17'd11355;
    value[8349] = 17'd11337;
    value[8350] = 17'd11320;
    value[8351] = 17'd11302;
    value[8352] = 17'd11285;
    value[8353] = 17'd11268;
    value[8354] = 17'd11250;
    value[8355] = 17'd11233;
    value[8356] = 17'd11216;
    value[8357] = 17'd11198;
    value[8358] = 17'd11181;
    value[8359] = 17'd11164;
    value[8360] = 17'd11146;
    value[8361] = 17'd11129;
    value[8362] = 17'd11112;
    value[8363] = 17'd11094;
    value[8364] = 17'd11077;
    value[8365] = 17'd11060;
    value[8366] = 17'd11042;
    value[8367] = 17'd11025;
    value[8368] = 17'd11008;
    value[8369] = 17'd10990;
    value[8370] = 17'd10973;
    value[8371] = 17'd10956;
    value[8372] = 17'd10938;
    value[8373] = 17'd10921;
    value[8374] = 17'd10904;
    value[8375] = 17'd10886;
    value[8376] = 17'd10869;
    value[8377] = 17'd10851;
    value[8378] = 17'd10834;
    value[8379] = 17'd10817;
    value[8380] = 17'd10799;
    value[8381] = 17'd10782;
    value[8382] = 17'd10765;
    value[8383] = 17'd10747;
    value[8384] = 17'd10730;
    value[8385] = 17'd10713;
    value[8386] = 17'd10695;
    value[8387] = 17'd10678;
    value[8388] = 17'd10661;
    value[8389] = 17'd10643;
    value[8390] = 17'd10626;
    value[8391] = 17'd10609;
    value[8392] = 17'd10591;
    value[8393] = 17'd10574;
    value[8394] = 17'd10556;
    value[8395] = 17'd10539;
    value[8396] = 17'd10522;
    value[8397] = 17'd10504;
    value[8398] = 17'd10487;
    value[8399] = 17'd10470;
    value[8400] = 17'd10452;
    value[8401] = 17'd10435;
    value[8402] = 17'd10418;
    value[8403] = 17'd10400;
    value[8404] = 17'd10383;
    value[8405] = 17'd10366;
    value[8406] = 17'd10348;
    value[8407] = 17'd10331;
    value[8408] = 17'd10313;
    value[8409] = 17'd10296;
    value[8410] = 17'd10279;
    value[8411] = 17'd10261;
    value[8412] = 17'd10244;
    value[8413] = 17'd10227;
    value[8414] = 17'd10209;
    value[8415] = 17'd10192;
    value[8416] = 17'd10175;
    value[8417] = 17'd10157;
    value[8418] = 17'd10140;
    value[8419] = 17'd10122;
    value[8420] = 17'd10105;
    value[8421] = 17'd10088;
    value[8422] = 17'd10070;
    value[8423] = 17'd10053;
    value[8424] = 17'd10036;
    value[8425] = 17'd10018;
    value[8426] = 17'd10001;
    value[8427] = 17'd09984;
    value[8428] = 17'd09966;
    value[8429] = 17'd09949;
    value[8430] = 17'd09931;
    value[8431] = 17'd09914;
    value[8432] = 17'd09897;
    value[8433] = 17'd09879;
    value[8434] = 17'd09862;
    value[8435] = 17'd09845;
    value[8436] = 17'd09827;
    value[8437] = 17'd09810;
    value[8438] = 17'd09793;
    value[8439] = 17'd09775;
    value[8440] = 17'd09758;
    value[8441] = 17'd09740;
    value[8442] = 17'd09723;
    value[8443] = 17'd09706;
    value[8444] = 17'd09688;
    value[8445] = 17'd09671;
    value[8446] = 17'd09654;
    value[8447] = 17'd09636;
    value[8448] = 17'd09619;
    value[8449] = 17'd09601;
    value[8450] = 17'd09584;
    value[8451] = 17'd09567;
    value[8452] = 17'd09549;
    value[8453] = 17'd09532;
    value[8454] = 17'd09515;
    value[8455] = 17'd09497;
    value[8456] = 17'd09480;
    value[8457] = 17'd09462;
    value[8458] = 17'd09445;
    value[8459] = 17'd09428;
    value[8460] = 17'd09410;
    value[8461] = 17'd09393;
    value[8462] = 17'd09376;
    value[8463] = 17'd09358;
    value[8464] = 17'd09341;
    value[8465] = 17'd09323;
    value[8466] = 17'd09306;
    value[8467] = 17'd09289;
    value[8468] = 17'd09271;
    value[8469] = 17'd09254;
    value[8470] = 17'd09237;
    value[8471] = 17'd09219;
    value[8472] = 17'd09202;
    value[8473] = 17'd09184;
    value[8474] = 17'd09167;
    value[8475] = 17'd09150;
    value[8476] = 17'd09132;
    value[8477] = 17'd09115;
    value[8478] = 17'd09098;
    value[8479] = 17'd09080;
    value[8480] = 17'd09063;
    value[8481] = 17'd09045;
    value[8482] = 17'd09028;
    value[8483] = 17'd09011;
    value[8484] = 17'd08993;
    value[8485] = 17'd08976;
    value[8486] = 17'd08958;
    value[8487] = 17'd08941;
    value[8488] = 17'd08924;
    value[8489] = 17'd08906;
    value[8490] = 17'd08889;
    value[8491] = 17'd08872;
    value[8492] = 17'd08854;
    value[8493] = 17'd08837;
    value[8494] = 17'd08819;
    value[8495] = 17'd08802;
    value[8496] = 17'd08785;
    value[8497] = 17'd08767;
    value[8498] = 17'd08750;
    value[8499] = 17'd08732;
    value[8500] = 17'd08715;
    value[8501] = 17'd08698;
    value[8502] = 17'd08680;
    value[8503] = 17'd08663;
    value[8504] = 17'd08646;
    value[8505] = 17'd08628;
    value[8506] = 17'd08611;
    value[8507] = 17'd08593;
    value[8508] = 17'd08576;
    value[8509] = 17'd08559;
    value[8510] = 17'd08541;
    value[8511] = 17'd08524;
    value[8512] = 17'd08506;
    value[8513] = 17'd08489;
    value[8514] = 17'd08472;
    value[8515] = 17'd08454;
    value[8516] = 17'd08437;
    value[8517] = 17'd08419;
    value[8518] = 17'd08402;
    value[8519] = 17'd08385;
    value[8520] = 17'd08367;
    value[8521] = 17'd08350;
    value[8522] = 17'd08333;
    value[8523] = 17'd08315;
    value[8524] = 17'd08298;
    value[8525] = 17'd08280;
    value[8526] = 17'd08263;
    value[8527] = 17'd08246;
    value[8528] = 17'd08228;
    value[8529] = 17'd08211;
    value[8530] = 17'd08193;
    value[8531] = 17'd08176;
    value[8532] = 17'd08159;
    value[8533] = 17'd08141;
    value[8534] = 17'd08124;
    value[8535] = 17'd08106;
    value[8536] = 17'd08089;
    value[8537] = 17'd08072;
    value[8538] = 17'd08054;
    value[8539] = 17'd08037;
    value[8540] = 17'd08019;
    value[8541] = 17'd08002;
    value[8542] = 17'd07985;
    value[8543] = 17'd07967;
    value[8544] = 17'd07950;
    value[8545] = 17'd07932;
    value[8546] = 17'd07915;
    value[8547] = 17'd07898;
    value[8548] = 17'd07880;
    value[8549] = 17'd07863;
    value[8550] = 17'd07845;
    value[8551] = 17'd07828;
    value[8552] = 17'd07811;
    value[8553] = 17'd07793;
    value[8554] = 17'd07776;
    value[8555] = 17'd07758;
    value[8556] = 17'd07741;
    value[8557] = 17'd07724;
    value[8558] = 17'd07706;
    value[8559] = 17'd07689;
    value[8560] = 17'd07671;
    value[8561] = 17'd07654;
    value[8562] = 17'd07637;
    value[8563] = 17'd07619;
    value[8564] = 17'd07602;
    value[8565] = 17'd07584;
    value[8566] = 17'd07567;
    value[8567] = 17'd07550;
    value[8568] = 17'd07532;
    value[8569] = 17'd07515;
    value[8570] = 17'd07497;
    value[8571] = 17'd07480;
    value[8572] = 17'd07463;
    value[8573] = 17'd07445;
    value[8574] = 17'd07428;
    value[8575] = 17'd07410;
    value[8576] = 17'd07393;
    value[8577] = 17'd07376;
    value[8578] = 17'd07358;
    value[8579] = 17'd07341;
    value[8580] = 17'd07323;
    value[8581] = 17'd07306;
    value[8582] = 17'd07289;
    value[8583] = 17'd07271;
    value[8584] = 17'd07254;
    value[8585] = 17'd07236;
    value[8586] = 17'd07219;
    value[8587] = 17'd07201;
    value[8588] = 17'd07184;
    value[8589] = 17'd07167;
    value[8590] = 17'd07149;
    value[8591] = 17'd07132;
    value[8592] = 17'd07114;
    value[8593] = 17'd07097;
    value[8594] = 17'd07080;
    value[8595] = 17'd07062;
    value[8596] = 17'd07045;
    value[8597] = 17'd07027;
    value[8598] = 17'd07010;
    value[8599] = 17'd06993;
    value[8600] = 17'd06975;
    value[8601] = 17'd06958;
    value[8602] = 17'd06940;
    value[8603] = 17'd06923;
    value[8604] = 17'd06906;
    value[8605] = 17'd06888;
    value[8606] = 17'd06871;
    value[8607] = 17'd06853;
    value[8608] = 17'd06836;
    value[8609] = 17'd06818;
    value[8610] = 17'd06801;
    value[8611] = 17'd06784;
    value[8612] = 17'd06766;
    value[8613] = 17'd06749;
    value[8614] = 17'd06731;
    value[8615] = 17'd06714;
    value[8616] = 17'd06697;
    value[8617] = 17'd06679;
    value[8618] = 17'd06662;
    value[8619] = 17'd06644;
    value[8620] = 17'd06627;
    value[8621] = 17'd06609;
    value[8622] = 17'd06592;
    value[8623] = 17'd06575;
    value[8624] = 17'd06557;
    value[8625] = 17'd06540;
    value[8626] = 17'd06522;
    value[8627] = 17'd06505;
    value[8628] = 17'd06488;
    value[8629] = 17'd06470;
    value[8630] = 17'd06453;
    value[8631] = 17'd06435;
    value[8632] = 17'd06418;
    value[8633] = 17'd06400;
    value[8634] = 17'd06383;
    value[8635] = 17'd06366;
    value[8636] = 17'd06348;
    value[8637] = 17'd06331;
    value[8638] = 17'd06313;
    value[8639] = 17'd06296;
    value[8640] = 17'd06279;
    value[8641] = 17'd06261;
    value[8642] = 17'd06244;
    value[8643] = 17'd06226;
    value[8644] = 17'd06209;
    value[8645] = 17'd06191;
    value[8646] = 17'd06174;
    value[8647] = 17'd06157;
    value[8648] = 17'd06139;
    value[8649] = 17'd06122;
    value[8650] = 17'd06104;
    value[8651] = 17'd06087;
    value[8652] = 17'd06070;
    value[8653] = 17'd06052;
    value[8654] = 17'd06035;
    value[8655] = 17'd06017;
    value[8656] = 17'd06000;
    value[8657] = 17'd05982;
    value[8658] = 17'd05965;
    value[8659] = 17'd05948;
    value[8660] = 17'd05930;
    value[8661] = 17'd05913;
    value[8662] = 17'd05895;
    value[8663] = 17'd05878;
    value[8664] = 17'd05860;
    value[8665] = 17'd05843;
    value[8666] = 17'd05826;
    value[8667] = 17'd05808;
    value[8668] = 17'd05791;
    value[8669] = 17'd05773;
    value[8670] = 17'd05756;
    value[8671] = 17'd05738;
    value[8672] = 17'd05721;
    value[8673] = 17'd05704;
    value[8674] = 17'd05686;
    value[8675] = 17'd05669;
    value[8676] = 17'd05651;
    value[8677] = 17'd05634;
    value[8678] = 17'd05617;
    value[8679] = 17'd05599;
    value[8680] = 17'd05582;
    value[8681] = 17'd05564;
    value[8682] = 17'd05547;
    value[8683] = 17'd05529;
    value[8684] = 17'd05512;
    value[8685] = 17'd05495;
    value[8686] = 17'd05477;
    value[8687] = 17'd05460;
    value[8688] = 17'd05442;
    value[8689] = 17'd05425;
    value[8690] = 17'd05407;
    value[8691] = 17'd05390;
    value[8692] = 17'd05373;
    value[8693] = 17'd05355;
    value[8694] = 17'd05338;
    value[8695] = 17'd05320;
    value[8696] = 17'd05303;
    value[8697] = 17'd05285;
    value[8698] = 17'd05268;
    value[8699] = 17'd05251;
    value[8700] = 17'd05233;
    value[8701] = 17'd05216;
    value[8702] = 17'd05198;
    value[8703] = 17'd05181;
    value[8704] = 17'd05163;
    value[8705] = 17'd05146;
    value[8706] = 17'd05129;
    value[8707] = 17'd05111;
    value[8708] = 17'd05094;
    value[8709] = 17'd05076;
    value[8710] = 17'd05059;
    value[8711] = 17'd05041;
    value[8712] = 17'd05024;
    value[8713] = 17'd05007;
    value[8714] = 17'd04989;
    value[8715] = 17'd04972;
    value[8716] = 17'd04954;
    value[8717] = 17'd04937;
    value[8718] = 17'd04919;
    value[8719] = 17'd04902;
    value[8720] = 17'd04884;
    value[8721] = 17'd04867;
    value[8722] = 17'd04850;
    value[8723] = 17'd04832;
    value[8724] = 17'd04815;
    value[8725] = 17'd04797;
    value[8726] = 17'd04780;
    value[8727] = 17'd04762;
    value[8728] = 17'd04745;
    value[8729] = 17'd04728;
    value[8730] = 17'd04710;
    value[8731] = 17'd04693;
    value[8732] = 17'd04675;
    value[8733] = 17'd04658;
    value[8734] = 17'd04640;
    value[8735] = 17'd04623;
    value[8736] = 17'd04606;
    value[8737] = 17'd04588;
    value[8738] = 17'd04571;
    value[8739] = 17'd04553;
    value[8740] = 17'd04536;
    value[8741] = 17'd04518;
    value[8742] = 17'd04501;
    value[8743] = 17'd04483;
    value[8744] = 17'd04466;
    value[8745] = 17'd04449;
    value[8746] = 17'd04431;
    value[8747] = 17'd04414;
    value[8748] = 17'd04396;
    value[8749] = 17'd04379;
    value[8750] = 17'd04361;
    value[8751] = 17'd04344;
    value[8752] = 17'd04327;
    value[8753] = 17'd04309;
    value[8754] = 17'd04292;
    value[8755] = 17'd04274;
    value[8756] = 17'd04257;
    value[8757] = 17'd04239;
    value[8758] = 17'd04222;
    value[8759] = 17'd04205;
    value[8760] = 17'd04187;
    value[8761] = 17'd04170;
    value[8762] = 17'd04152;
    value[8763] = 17'd04135;
    value[8764] = 17'd04117;
    value[8765] = 17'd04100;
    value[8766] = 17'd04082;
    value[8767] = 17'd04065;
    value[8768] = 17'd04048;
    value[8769] = 17'd04030;
    value[8770] = 17'd04013;
    value[8771] = 17'd03995;
    value[8772] = 17'd03978;
    value[8773] = 17'd03960;
    value[8774] = 17'd03943;
    value[8775] = 17'd03925;
    value[8776] = 17'd03908;
    value[8777] = 17'd03891;
    value[8778] = 17'd03873;
    value[8779] = 17'd03856;
    value[8780] = 17'd03838;
    value[8781] = 17'd03821;
    value[8782] = 17'd03803;
    value[8783] = 17'd03786;
    value[8784] = 17'd03769;
    value[8785] = 17'd03751;
    value[8786] = 17'd03734;
    value[8787] = 17'd03716;
    value[8788] = 17'd03699;
    value[8789] = 17'd03681;
    value[8790] = 17'd03664;
    value[8791] = 17'd03646;
    value[8792] = 17'd03629;
    value[8793] = 17'd03612;
    value[8794] = 17'd03594;
    value[8795] = 17'd03577;
    value[8796] = 17'd03559;
    value[8797] = 17'd03542;
    value[8798] = 17'd03524;
    value[8799] = 17'd03507;
    value[8800] = 17'd03489;
    value[8801] = 17'd03472;
    value[8802] = 17'd03455;
    value[8803] = 17'd03437;
    value[8804] = 17'd03420;
    value[8805] = 17'd03402;
    value[8806] = 17'd03385;
    value[8807] = 17'd03367;
    value[8808] = 17'd03350;
    value[8809] = 17'd03332;
    value[8810] = 17'd03315;
    value[8811] = 17'd03298;
    value[8812] = 17'd03280;
    value[8813] = 17'd03263;
    value[8814] = 17'd03245;
    value[8815] = 17'd03228;
    value[8816] = 17'd03210;
    value[8817] = 17'd03193;
    value[8818] = 17'd03175;
    value[8819] = 17'd03158;
    value[8820] = 17'd03141;
    value[8821] = 17'd03123;
    value[8822] = 17'd03106;
    value[8823] = 17'd03088;
    value[8824] = 17'd03071;
    value[8825] = 17'd03053;
    value[8826] = 17'd03036;
    value[8827] = 17'd03018;
    value[8828] = 17'd03001;
    value[8829] = 17'd02984;
    value[8830] = 17'd02966;
    value[8831] = 17'd02949;
    value[8832] = 17'd02931;
    value[8833] = 17'd02914;
    value[8834] = 17'd02896;
    value[8835] = 17'd02879;
    value[8836] = 17'd02861;
    value[8837] = 17'd02844;
    value[8838] = 17'd02827;
    value[8839] = 17'd02809;
    value[8840] = 17'd02792;
    value[8841] = 17'd02774;
    value[8842] = 17'd02757;
    value[8843] = 17'd02739;
    value[8844] = 17'd02722;
    value[8845] = 17'd02704;
    value[8846] = 17'd02687;
    value[8847] = 17'd02670;
    value[8848] = 17'd02652;
    value[8849] = 17'd02635;
    value[8850] = 17'd02617;
    value[8851] = 17'd02600;
    value[8852] = 17'd02582;
    value[8853] = 17'd02565;
    value[8854] = 17'd02547;
    value[8855] = 17'd02530;
    value[8856] = 17'd02513;
    value[8857] = 17'd02495;
    value[8858] = 17'd02478;
    value[8859] = 17'd02460;
    value[8860] = 17'd02443;
    value[8861] = 17'd02425;
    value[8862] = 17'd02408;
    value[8863] = 17'd02390;
    value[8864] = 17'd02373;
    value[8865] = 17'd02355;
    value[8866] = 17'd02338;
    value[8867] = 17'd02321;
    value[8868] = 17'd02303;
    value[8869] = 17'd02286;
    value[8870] = 17'd02268;
    value[8871] = 17'd02251;
    value[8872] = 17'd02233;
    value[8873] = 17'd02216;
    value[8874] = 17'd02198;
    value[8875] = 17'd02181;
    value[8876] = 17'd02164;
    value[8877] = 17'd02146;
    value[8878] = 17'd02129;
    value[8879] = 17'd02111;
    value[8880] = 17'd02094;
    value[8881] = 17'd02076;
    value[8882] = 17'd02059;
    value[8883] = 17'd02041;
    value[8884] = 17'd02024;
    value[8885] = 17'd02006;
    value[8886] = 17'd01989;
    value[8887] = 17'd01972;
    value[8888] = 17'd01954;
    value[8889] = 17'd01937;
    value[8890] = 17'd01919;
    value[8891] = 17'd01902;
    value[8892] = 17'd01884;
    value[8893] = 17'd01867;
    value[8894] = 17'd01849;
    value[8895] = 17'd01832;
    value[8896] = 17'd01815;
    value[8897] = 17'd01797;
    value[8898] = 17'd01780;
    value[8899] = 17'd01762;
    value[8900] = 17'd01745;
    value[8901] = 17'd01727;
    value[8902] = 17'd01710;
    value[8903] = 17'd01692;
    value[8904] = 17'd01675;
    value[8905] = 17'd01657;
    value[8906] = 17'd01640;
    value[8907] = 17'd01623;
    value[8908] = 17'd01605;
    value[8909] = 17'd01588;
    value[8910] = 17'd01570;
    value[8911] = 17'd01553;
    value[8912] = 17'd01535;
    value[8913] = 17'd01518;
    value[8914] = 17'd01500;
    value[8915] = 17'd01483;
    value[8916] = 17'd01466;
    value[8917] = 17'd01448;
    value[8918] = 17'd01431;
    value[8919] = 17'd01413;
    value[8920] = 17'd01396;
    value[8921] = 17'd01378;
    value[8922] = 17'd01361;
    value[8923] = 17'd01343;
    value[8924] = 17'd01326;
    value[8925] = 17'd01308;
    value[8926] = 17'd01291;
    value[8927] = 17'd01274;
    value[8928] = 17'd01256;
    value[8929] = 17'd01239;
    value[8930] = 17'd01221;
    value[8931] = 17'd01204;
    value[8932] = 17'd01186;
    value[8933] = 17'd01169;
    value[8934] = 17'd01151;
    value[8935] = 17'd01134;
    value[8936] = 17'd01116;
    value[8937] = 17'd01099;
    value[8938] = 17'd01082;
    value[8939] = 17'd01064;
    value[8940] = 17'd01047;
    value[8941] = 17'd01029;
    value[8942] = 17'd01012;
    value[8943] = 17'd00994;
    value[8944] = 17'd00977;
    value[8945] = 17'd00959;
    value[8946] = 17'd00942;
    value[8947] = 17'd00925;
    value[8948] = 17'd00907;
    value[8949] = 17'd00890;
    value[8950] = 17'd00872;
    value[8951] = 17'd00855;
    value[8952] = 17'd00837;
    value[8953] = 17'd00820;
    value[8954] = 17'd00802;
    value[8955] = 17'd00785;
    value[8956] = 17'd00767;
    value[8957] = 17'd00750;
    value[8958] = 17'd00733;
    value[8959] = 17'd00715;
    value[8960] = 17'd00698;
    value[8961] = 17'd00680;
    value[8962] = 17'd00663;
    value[8963] = 17'd00645;
    value[8964] = 17'd00628;
    value[8965] = 17'd00610;
    value[8966] = 17'd00593;
    value[8967] = 17'd00575;
    value[8968] = 17'd00558;
    value[8969] = 17'd00541;
    value[8970] = 17'd00523;
    value[8971] = 17'd00506;
    value[8972] = 17'd00488;
    value[8973] = 17'd00471;
    value[8974] = 17'd00453;
    value[8975] = 17'd00436;
    value[8976] = 17'd00418;
    value[8977] = 17'd00401;
    value[8978] = 17'd00383;
    value[8979] = 17'd00366;
    value[8980] = 17'd00349;
    value[8981] = 17'd00331;
    value[8982] = 17'd00314;
    value[8983] = 17'd00296;
    value[8984] = 17'd00279;
    value[8985] = 17'd00261;
    value[8986] = 17'd00244;
    value[8987] = 17'd00226;
    value[8988] = 17'd00209;
    value[8989] = 17'd00191;
    value[8990] = 17'd00174;
    value[8991] = 17'd00157;
    value[8992] = 17'd00139;
    value[8993] = 17'd00122;
    value[8994] = 17'd00104;
    value[8995] = 17'd00087;
    value[8996] = 17'd00069;
    value[8997] = 17'd00052;
    value[8998] = 17'd00034;
    value[8999] = 17'd00017;
    value[9000] = 17'd00000;
  end

endmodule
